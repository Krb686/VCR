library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity SAMPLE_PLAYBACK is
    Port ( clk : in  STD_LOGIC;
           rst : in  STD_LOGIC;
           dout : out  STD_LOGIC_VECTOR (11 downto 0));
end SAMPLE_PLAYBACK;

architecture Behavioral of SAMPLE_PLAYBACK is

	--constant ROM_LENGTH	: integer	:= 576;				-- small blip
	--constant ROM_LENGTH	: integer	:= 4096;			-- open
	constant ROM_LENGTH	:	integer	:= 4656;				-- up_2

	type ROM is array (0 to ROM_LENGTH - 1) of std_logic_vector(11 downto 0);
	
--				constant DATA_ROM	: ROM := ( 
--			x"3c9", x"3c5", x"3bf", x"3bf", x"3c2", x"3ba", x"3af", x"3ae", x"3b6", x"3af", x"3b2", x"3b2", x"45e", x"3aa", x"45e", x"3b8", 
--			x"4de", x"38e", x"438", x"385", x"39a", x"3ab", x"464", x"39d", x"390", x"396", x"448", x"4f2", x"397", x"386", x"38b", x"39e", 
--			x"4b1", x"3c3", x"3b2", x"3a2", x"38d", x"39d", x"3a0", x"3a9", x"39c", x"39b", x"258", x"3a5", x"3a1", x"3b0", x"3b7", x"271",  --first sample to be loaded is 3b0
--			x"3b8", x"3c6", x"3c4", x"3c7", x"3be", x"3bd", x"3bf", x"3c9", x"3d6", x"3de", x"3de", x"3d4", x"3df", x"3ec", x"3f2", x"3f8", 
--			x"3f5", x"3ec", x"3de", x"3de", x"3df", x"3f4", x"3ed", x"3e5", x"3d3", x"3cb", x"3c1", x"3c7", x"3cc", x"3c3", x"3bd", x"3af", 
--			x"3ad", x"3a6", x"3a6", x"39d", x"3a0", x"391", x"38d", x"37b", x"372", x"36d", x"361", x"35e", x"356", x"343", x"334", x"329", 
--			x"323", x"31f", x"321", x"320", x"323", x"31e", x"317", x"303", x"2f9", x"2f6", x"30b", x"334", x"368", x"39c", x"3ef", x"424", 
--			x"44d", x"466", x"463", x"44f", x"442", x"438", x"42d", x"433", x"438", x"448", x"448", x"45b", x"45e", x"464", x"463", x"459", 
--			x"44e", x"444", x"434", x"427", x"418", x"40b", x"405", x"3fd", x"3f2", x"3e5", x"3d9", x"3c8", x"3ba", x"3aa", x"39f", x"38b", 
--			x"375", x"362", x"34b", x"335", x"321", x"316", x"2fb", x"2e4", x"2cf", x"2c6", x"2c8", x"2c7", x"2c9", x"2c4", x"2c1", x"2e4", 
--			x"332", x"3ea", x"463", x"4cc", x"4ad", x"46a", x"3f9", x"3e2", x"3c8", x"3dd", x"3e4", x"3dc", x"3a4", x"396", x"39c", x"3aa", 
--			x"3f0", x"407", x"420", x"404", x"3f8", x"3cd", x"3dc", x"3e1", x"3f6", x"3de", x"3cf", x"3a2", x"390", x"38d", x"3ac", x"3fc",
--			x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac",
--			x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac",
--			x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac",
--			x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac",
--			x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac",
--			x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac",
--			x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac",
--			x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac",
--			x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac",
--			x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac",
--			x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac",
--			x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac",
--			x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac",
--			x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac",
--			x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac",
--			x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac",
--			x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac",
--			x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac",
--			x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac",
--			x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac",
--			x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac",
--			x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac",
--			x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac",
--			x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac", x"3ac" 			
--			);





--				constant DATA_ROM : ROM := ( 
--			x"3aa", x"3af", x"3ab", x"3ab", x"3ad", x"3a8", x"3aa", x"3aa", x"3ab", x"3ba", x"3ab", x"3a9", x"39c", x"39e", x"39e", x"39f", 
--			x"39d", x"38c", x"391", x"396", x"3a6", x"3af", x"3b3", x"39c", x"394", x"394", x"3a3", x"3a4", x"3a5", x"3a7", x"3ab", x"3a5", 
--			x"3a6", x"39f", x"39d", x"39d", x"3a7", x"39d", x"3ad", x"3ae", x"3b3", x"3a9", x"3ac", x"3af", x"3b9", x"3b8", x"3a6", x"393", 
--			x"386", x"39e", x"3b6", x"3c7", x"3cb", x"3be", x"3be", x"3b4", x"3b6", x"3ad", x"3b2", x"3af", x"3b6", x"3c3", x"3d0", x"3da", 
--			x"3c9", x"3c5", x"3bf", x"3bf", x"3c2", x"3ba", x"3af", x"3ae", x"3b6", x"3af", x"3b2", x"3b2", x"3ab", x"3aa", x"3b2", x"3b8", 
--			x"3a4", x"38e", x"38b", x"385", x"39a", x"3ab", x"3a8", x"39d", x"390", x"396", x"3a1", x"3a4", x"397", x"386", x"38b", x"39e", 
--			x"3ac", x"3c3", x"3b2", x"3a2", x"38d", x"39d", x"3a0", x"3a9", x"39c", x"39b", x"3a2", x"3a5", x"3a1", x"3b0", x"3b7", x"3ab", 
--			x"3b8", x"3c6", x"3c4", x"3c7", x"3be", x"3bd", x"3bf", x"3c9", x"3d6", x"3de", x"3de", x"3d4", x"3df", x"3ec", x"3f2", x"3f8", 
--			x"3f5", x"3ec", x"3de", x"3de", x"3df", x"3f4", x"3ed", x"3e5", x"3d3", x"3cb", x"3c1", x"3c7", x"3cc", x"3c3", x"3bd", x"3af", 
--			x"3ad", x"3a6", x"3a6", x"39d", x"3a0", x"391", x"38d", x"37b", x"372", x"36d", x"361", x"35e", x"356", x"343", x"334", x"329", 
--			x"323", x"31f", x"321", x"320", x"323", x"31e", x"317", x"303", x"2f9", x"2f6", x"30b", x"334", x"368", x"39c", x"3ef", x"424", 
--			x"44d", x"466", x"463", x"44f", x"442", x"438", x"42d", x"433", x"438", x"448", x"448", x"45b", x"45e", x"464", x"463", x"459", 
--			x"44e", x"444", x"434", x"427", x"418", x"40b", x"405", x"3fd", x"3f2", x"3e5", x"3d9", x"3c8", x"3ba", x"3aa", x"39f", x"38b", 
--			x"375", x"362", x"34b", x"335", x"321", x"316", x"2fb", x"2e4", x"2cf", x"2c6", x"2c8", x"2c7", x"2c9", x"2c4", x"2c1", x"2e4", 
--			x"332", x"3ea", x"463", x"4cc", x"4ad", x"46a", x"3f9", x"3e2", x"3c8", x"3dd", x"3e4", x"3dc", x"3a4", x"396", x"39c", x"3aa", 
--			x"3f0", x"407", x"420", x"404", x"3f8", x"3cd", x"3dc", x"3e1", x"3f6", x"3de", x"3cf", x"3a2", x"390", x"38d", x"3ac", x"3fc", 
--			x"429", x"43c", x"41a", x"3fd", x"3d2", x"3e8", x"3f5", x"40e", x"40c", x"3fd", x"3d3", x"3cd", x"3cb", x"3db", x"3e5", x"3e5", 
--			x"3c5", x"3ab", x"397", x"384", x"388", x"383", x"370", x"356", x"337", x"30c", x"2f8", x"2e1", x"2da", x"2da", x"2da", x"2cf", 
--			x"2c6", x"2db", x"306", x"370", x"40b", x"46c", x"4b8", x"4a5", x"46f", x"41e", x"40c", x"3e7", x"3ee", x"3e4", x"3d0", x"392", 
--			x"372", x"34d", x"352", x"371", x"39d", x"3c1", x"3df", x"3de", x"3d4", x"3dc", x"3de", x"3f9", x"3fd", x"3fd", x"3d2", x"3b2", 
--			x"387", x"37f", x"386", x"3c0", x"3f0", x"422", x"42b", x"41c", x"40a", x"3f7", x"404", x"40b", x"420", x"418", x"40d", x"3eb", 
--			x"3cf", x"3b2", x"3a5", x"39e", x"39f", x"38d", x"38a", x"373", x"362", x"359", x"34e", x"348", x"333", x"311", x"2ec", x"2cb", 
--			x"2b3", x"2a8", x"2a3", x"2b5", x"2d8", x"33b", x"3b5", x"42a", x"499", x"4b3", x"4a7", x"46f", x"456", x"422", x"421", x"404", 
--			x"3f6", x"3ac", x"37f", x"338", x"31e", x"31e", x"333", x"35e", x"38d", x"3ae", x"3bf", x"3d9", x"3e2", x"406", x"41a", x"433", 
--			x"423", x"411", x"3da", x"3b1", x"38a", x"37f", x"388", x"3a8", x"3cb", x"3e8", x"3fb", x"3f6", x"3f8", x"401", x"40a", x"423", 
--			x"433", x"42d", x"41c", x"3f8", x"3cd", x"3a4", x"394", x"386", x"379", x"37a", x"368", x"35c", x"350", x"33e", x"340", x"341", 
--			x"335", x"327", x"309", x"2e4", x"2c3", x"2a4", x"2ae", x"2d1", x"331", x"39e", x"409", x"468", x"47f", x"482", x"462", x"454", 
--			x"43c", x"448", x"436", x"426", x"3e1", x"3a4", x"355", x"325", x"311", x"31c", x"33d", x"35c", x"380", x"396", x"3b5", x"3bf", 
--			x"3e8", x"40e", x"430", x"43d", x"43d", x"41b", x"3f1", x"3bd", x"39e", x"397", x"39a", x"3ac", x"3b7", x"3cc", x"3ca", x"3d7", 
--			x"3d8", x"3e9", x"409", x"424", x"434", x"439", x"41d", x"3fe", x"3d6", x"3b0", x"39c", x"38a", x"380", x"372", x"35f", x"34b", 
--			x"33b", x"331", x"336", x"32e", x"32b", x"315", x"2fa", x"2db", x"2ba", x"2b3", x"2ca", x"31b", x"379", x"3e9", x"447", x"46c", 
--			x"473", x"454", x"44b", x"430", x"44a", x"43f", x"43d", x"412", x"3d8", x"381", x"348", x"31a", x"311", x"324", x"34a", x"368", 
--			x"385", x"39c", x"3a5", x"3c7", x"3df", x"40e", x"42e", x"445", x"43c", x"42a", x"3fe", x"3cd", x"3a3", x"38d", x"38a", x"390", 
--			x"3a9", x"3b7", x"3c1", x"3c4", x"3d5", x"3e7", x"409", x"422", x"438", x"437", x"42e", x"409", x"3ea", x"3c6", x"3ac", x"39f", 
--			x"38d", x"381", x"370", x"35f", x"349", x"341", x"344", x"34f", x"349", x"344", x"32a", x"30d", x"2e6", x"2c4", x"2b7", x"2c1", 
--			x"30b", x"359", x"3bf", x"41b", x"449", x"45a", x"450", x"443", x"435", x"44c", x"452", x"457", x"437", x"401", x"3b1", x"371", 
--			x"331", x"31e", x"31e", x"332", x"34d", x"368", x"381", x"38a", x"3a4", x"3b5", x"3e1", x"405", x"430", x"43b", x"43d", x"421", 
--			x"3fe", x"3d5", x"3ac", x"394", x"397", x"39f", x"3b0", x"3bf", x"3c1", x"3cb", x"3d3", x"3e1", x"3f1", x"412", x"41f", x"426", 
--			x"41b", x"402", x"3e8", x"3ce", x"3b3", x"3a8", x"398", x"38a", x"37b", x"362", x"356", x"343", x"33d", x"33e", x"335", x"32b", 
--			x"311", x"2f7", x"2d5", x"2b5", x"2b1", x"2d5", x"31d", x"36d", x"3d5", x"41d", x"44d", x"44a", x"449", x"43c", x"442", x"44d", 
--			x"453", x"456", x"435", x"3ff", x"3ad", x"36e", x"332", x"31d", x"31a", x"329", x"346", x"366", x"379", x"38d", x"398", x"3b4", 
--			x"3cd", x"3ec", x"413", x"424", x"435", x"422", x"40b", x"3e1", x"3c0", x"3a9", x"3aa", x"3af", x"3c3", x"3d2", x"3d8", x"3d6", 
--			x"3d0", x"3d1", x"3df", x"3ef", x"400", x"414", x"40f", x"405", x"3f0", x"3cf", x"3b8", x"3a7", x"39f", x"399", x"387", x"377", 
--			x"361", x"350", x"342", x"338", x"330", x"322", x"310", x"2fa", x"2df", x"2c2", x"2b9", x"2ca", x"2fd", x"344", x"3a3", x"3fc", 
--			x"434", x"44e", x"44b", x"441", x"43c", x"448", x"448", x"455", x"444", x"422", x"3e3", x"39f", x"35d", x"332", x"321", x"322", 
--			x"339", x"356", x"36a", x"377", x"389", x"392", x"3a1", x"3bc", x"3e2", x"3fd", x"41b", x"424", x"420", x"409", x"3ea", x"3d5", 
--			x"3c8", x"3c8", x"3d4", x"3e2", x"3de", x"3da", x"3cb", x"3c2", x"3c5", x"3d2", x"3e5", x"3fa", x"404", x"403", x"3f6", x"3e2", 
--			x"3ca", x"3b9", x"3ad", x"3a4", x"3a5", x"392", x"380", x"36d", x"352", x"340", x"32f", x"324", x"31b", x"309", x"2f4", x"2db", 
--			x"2c3", x"2b5", x"2c8", x"2ff", x"33e", x"39c", x"3ed", x"425", x"43e", x"446", x"43a", x"437", x"444", x"44c", x"456", x"449", 
--			x"42e", x"3f9", x"3b9", x"378", x"34d", x"333", x"32f", x"336", x"349", x"355", x"366", x"36d", x"376", x"381", x"399", x"3ba", 
--			x"3dc", x"406", x"41b", x"423", x"415", x"40a", x"3f5", x"3e5", x"3e0", x"3e2", x"3e8", x"3e7", x"3e0", x"3d2", x"3ca", x"3c3", 
--			x"3c4", x"3d1", x"3df", x"3f0", x"3f7", x"3f1", x"3e0", x"3d4", x"3c7", x"3be", x"3b5", x"3ae", x"3a4", x"392", x"379", x"367", 
--			x"34f", x"340", x"332", x"328", x"316", x"30a", x"2f1", x"2da", x"2c3", x"2b5", x"2cd", x"2fc", x"33e", x"392", x"3da", x"411", 
--			x"42b", x"435", x"434", x"43b", x"445", x"453", x"45f", x"459", x"43d", x"40d", x"3d2", x"390", x"365", x"342", x"334", x"33a", 
--			x"340", x"347", x"356", x"35d", x"365", x"379", x"392", x"3af", x"3d2", x"3f7", x"412", x"41c", x"41f", x"413", x"40b", x"401", 
--			x"400", x"403", x"3ff", x"3f6", x"3e5", x"3d7", x"3cb", x"3bf", x"3c0", x"3cd", x"3d6", x"3df", x"3dd", x"3da", x"3d2", x"3c9", 
--			x"3c2", x"3b7", x"3b3", x"3a9", x"39e", x"397", x"37e", x"368", x"355", x"344", x"331", x"321", x"30b", x"2ef", x"2d1", x"2b8", 
--			x"2a5", x"2ae", x"2da", x"30f", x"366", x"3b2", x"3f4", x"420", x"434", x"43d", x"43d", x"44f", x"459", x"470", x"46b", x"459", 
--			x"42e", x"3f6", x"3b0", x"377", x"34a", x"333", x"331", x"339", x"341", x"353", x"35b", x"362", x"36e", x"379", x"394", x"3af", 
--			x"3da", x"3fb", x"416", x"420", x"422", x"41a", x"410", x"410", x"40a", x"40b", x"402", x"3fd", x"3e8", x"3de", x"3cf", x"3c9", 
--			x"3cc", x"3cc", x"3d5", x"3d9", x"3d7", x"3cc", x"3c2", x"3b3", x"3ae", x"3a9", x"3ad", x"3ac", x"3a4", x"39b", x"381", x"36e", 
--			x"34f", x"333", x"31a", x"2fd", x"2e6", x"2c9", x"2b2", x"29e", x"2a6", x"2d2", x"303", x"35c", x"3a3", x"3ee", x"41b", x"437", 
--			x"442", x"448", x"45f", x"461", x"475", x"474", x"462", x"435", x"3ff", x"3b9", x"37e", x"353", x"33b", x"338", x"33f", x"345", 
--			x"354", x"357", x"362", x"366", x"376", x"389", x"3a5", x"3d0", x"3f6", x"414", x"41d", x"420", x"41f", x"418", x"415", x"419", 
--			x"41a", x"410", x"40c", x"3fb", x"3ea", x"3d9", x"3cd", x"3cd", x"3cd", x"3d0", x"3d0", x"3ca", x"3c0", x"3b3", x"3ad", x"3ab", 
--			x"3ad", x"3ae", x"3ad", x"3a1", x"394", x"37f", x"366", x"34a", x"32c", x"30f", x"2f0", x"2d3", x"2af", x"295", x"285", x"2ad", 
--			x"2d4", x"31c", x"378", x"3bb", x"406", x"427", x"442", x"448", x"459", x"466", x"476", x"489", x"479", x"467", x"42b", x"3ec", 
--			x"3a9", x"372", x"34f", x"33a", x"33b", x"33b", x"34a", x"351", x"34a", x"354", x"35a", x"375", x"38d", x"3c4", x"3f2", x"419", 
--			x"42d", x"431", x"432", x"42b", x"426", x"422", x"428", x"417", x"411", x"3fa", x"3de", x"3cc", x"3bf", x"3ca", x"3d8", x"3dd", 
--			x"3e4", x"3e0", x"3d3", x"3c4", x"3c2", x"3ba", x"3c3", x"3bc", x"3bc", x"3a8", x"38d", x"36c", x"340", x"320", x"2f6", x"2d5", 
--			x"2af", x"286", x"263", x"246", x"246", x"298", x"2ed", x"36d", x"41f", x"48a", x"4c7", x"4ce", x"4b1", x"481", x"460", x"46e", 
--			x"44d", x"458", x"415", x"3c9", x"35a", x"2fe", x"2b8", x"2a9", x"2dc", x"30f", x"375", x"3a8", x"3de", x"3ea", x"3f3", x"403", 
--			x"41c", x"450", x"462", x"46d", x"445", x"3fb", x"3a3", x"354", x"33a", x"349", x"37a", x"3bb", x"3fc", x"40f", x"417", x"40b", 
--			x"405", x"430", x"456", x"47f", x"489", x"464", x"418", x"3c7", x"37c", x"35a", x"362", x"36d", x"37d", x"378", x"362", x"33f", 
--			x"331", x"33a", x"342", x"356", x"341", x"314", x"2cf", x"26c", x"231", x"219", x"24d", x"2f4", x"3a5", x"458", x"4e9", x"4e1", 
--			x"4c9", x"47c", x"453", x"433", x"443", x"43d", x"3ee", x"3a5", x"310", x"2bc", x"284", x"2ba", x"307", x"391", x"3f9", x"421", 
--			x"444", x"41e", x"425", x"42b", x"44d", x"455", x"43f", x"3f2", x"37a", x"32b", x"2e3", x"2e7", x"316", x"35c", x"39a", x"3f3", 
--			x"429", x"447", x"48a", x"480", x"499", x"485", x"462", x"42f", x"3f8", x"3bd", x"397", x"39c", x"38d", x"3a1", x"39d", x"39b", 
--			x"39e", x"3a3", x"3b1", x"3c4", x"3d5", x"3bf", x"3ae", x"37b", x"33d", x"302", x"2b8", x"281", x"246", x"222", x"201", x"214", 
--			x"263", x"340", x"41e", x"4e5", x"586", x"549", x"50c", x"47b", x"436", x"3e7", x"3e1", x"3b3", x"350", x"307", x"279", x"271", 
--			x"28a", x"328", x"3a1", x"449", x"49d", x"48a", x"485", x"441", x"441", x"42b", x"429", x"3e9", x"395", x"335", x"2c7", x"2c7", 
--			x"2d6", x"32e", x"386", x"3dc", x"41b", x"457", x"491", x"4a0", x"4c9", x"499", x"469", x"418", x"3c7", x"395", x"381", x"397", 
--			x"3aa", x"3c8", x"3bd", x"3b7", x"3b4", x"3b8", x"3d6", x"3ef", x"3f8", x"3d7", x"3b7", x"372", x"341", x"31f", x"2ed", x"2cb", 
--			x"285", x"25e", x"22b", x"21f", x"23b", x"279", x"343", x"433", x"4c8", x"567", x"53f", x"4ef", x"47b", x"42a", x"3e5", x"3ab", 
--			x"3a6", x"313", x"2e5", x"27e", x"27d", x"2bc", x"359", x"3f6", x"464", x"4c0", x"488", x"47c", x"452", x"43c", x"426", x"3f9", 
--			x"3a0", x"32a", x"2e9", x"2a9", x"2d0", x"323", x"379", x"3d6", x"407", x"444", x"480", x"4c8", x"4d4", x"4c4", x"471", x"3fb", 
--			x"3a2", x"378", x"388", x"3af", x"3d2", x"3d9", x"3d2", x"3bd", x"3c2", x"3df", x"405", x"41b", x"409", x"3df", x"393", x"36b", 
--			x"34b", x"338", x"326", x"2e2", x"2a6", x"261", x"230", x"225", x"23e", x"278", x"2bc", x"3b5", x"47d", x"42e", x"44d", x"452", 
--			x"448", x"412", x"3cd", x"38a", x"35d", x"35f", x"363", x"377", x"379", x"362", x"33d", x"30c", x"2e6", x"2c6", x"2c2", x"2f2", 
--			x"351", x"3b6", x"40e", x"43a", x"43a", x"415", x"3f7", x"3e2", x"3dc", x"3fe", x"41a", x"429", x"423", x"401", x"3de", x"3bb", 
--			x"3b9", x"3c1", x"3df", x"3fe", x"409", x"40b", x"3fd", x"3e9", x"3df", x"3de", x"3df", x"3e4", x"3e4", x"3d5", x"3be", x"3ae", 
--			x"3aa", x"3bd", x"3e0", x"3fe", x"409", x"408", x"3f9", x"3da", x"3c5", x"3be", x"3ca", x"3e4", x"3f6", x"3f7", x"3d7", x"3ac", 
--			x"380", x"35e", x"35a", x"357", x"364", x"358", x"337", x"309", x"2d4", x"2af", x"29a", x"2ae", x"2ed", x"33e", x"38f", x"3cb", 
--			x"3df", x"3d0", x"3af", x"39d", x"38e", x"39f", x"3c4", x"3dc", x"3ea", x"3dd", x"3bb", x"39c", x"387", x"390", x"39d", x"3c6", 
--			x"3e2", x"3f2", x"3ef", x"3d9", x"3be", x"39e", x"396", x"390", x"38e", x"395", x"38a", x"38e", x"38a", x"398", x"3a1", x"3aa", 
--			x"3b1", x"3b2", x"3b8", x"3b1", x"3b0", x"3b8", x"3b5", x"3b7", x"3a6", x"38d", x"370", x"351", x"341", x"334", x"33c", x"33b", 
--			x"337", x"32f", x"311", x"2f1", x"2da", x"2c9", x"2cc", x"2eb", x"31a", x"345", x"378", x"385", x"387", x"378", x"366", x"35a", 
--			x"35b", x"379", x"39a", x"3bd", x"3cf", x"3ce", x"3c2", x"3ac", x"3a1", x"39f", x"3aa", x"3c0", x"3d6", x"3d9", x"3cc", x"3ba", 
--			x"39a", x"382", x"37b", x"375", x"383", x"394", x"3aa", x"3ad", x"3b0", x"3a9", x"39e", x"395", x"38e", x"394", x"39b", x"39b", 
--			x"3a8", x"3a4", x"39f", x"389", x"379", x"369", x"35d", x"360", x"35a", x"354", x"34a", x"335", x"319", x"2f8", x"2db", x"2d0", 
--			x"2d1", x"2e4", x"306", x"332", x"353", x"36c", x"37a", x"37b", x"379", x"378", x"38a", x"393", x"3a9", x"3b7", x"3be", x"3b9", 
--			x"3aa", x"39d", x"392", x"38f", x"38e", x"398", x"3a1", x"3a6", x"3a9", x"39d", x"395", x"387", x"374", x"36a", x"368", x"36e", 
--			x"378", x"382", x"381", x"383", x"37d", x"376", x"379", x"377", x"389", x"39c", x"3b6", x"3c3", x"3c6", x"3ba", x"39e", x"38b", 
--			x"373", x"367", x"358", x"34f", x"344", x"321", x"2f9", x"2c6", x"29b", x"27d", x"267", x"264", x"268", x"272", x"288", x"292", 
--			x"29d", x"29c", x"2a2", x"2ad", x"2c3", x"2de", x"2fb", x"322", x"346", x"364", x"37e", x"387", x"397", x"3a8", x"3c2", x"3dd", 
--			x"3f8", x"414", x"42c", x"438", x"43a", x"435", x"42f", x"425", x"422", x"423", x"423", x"42b", x"433", x"434", x"436", x"430", 
--			x"420", x"415", x"411", x"40a", x"406", x"3ff", x"3ee", x"3e1", x"3c6", x"3ba", x"3b1", x"3b1", x"3b8", x"3c0", x"3be", x"3b6", 
--			x"3a6", x"38f", x"36a", x"348", x"316", x"2ed", x"2b9", x"290", x"279", x"27c", x"28c", x"28a", x"28b", x"28d", x"29c", x"2b2", 
--			x"2d0", x"2fb", x"324", x"34e", x"36f", x"38e", x"3a1", x"3b0", x"3b7", x"3c4", x"3d2", x"3de", x"3ef", x"3fe", x"40c", x"40e", 
--			x"40d", x"40e", x"408", x"404", x"404", x"41a", x"424", x"42b", x"42a", x"41f", x"40d", x"404", x"3f7", x"3f2", x"3f8", x"3fc", 
--			x"3f9", x"3f1", x"3dc", x"3cb", x"3b1", x"39d", x"392", x"381", x"371", x"359", x"34a", x"334", x"31e", x"303", x"2e0", x"2bd", 
--			x"29e", x"286", x"288", x"29d", x"2c8", x"2ed", x"315", x"336", x"345", x"354", x"35c", x"361", x"361", x"370", x"374", x"378", 
--			x"37a", x"372", x"37b", x"389", x"39c", x"3ae", x"3ba", x"3c4", x"3c2", x"3b7", x"3aa", x"39a", x"388", x"37a", x"36a", x"366", 
--			x"36b", x"379", x"38c", x"39d", x"3a9", x"3b2", x"3be", x"3c4", x"3c9", x"3d4", x"3d9", x"3dc", x"3d9", x"3ce", x"3b9", x"3a9", 
--			x"39e", x"39b", x"3a6", x"3b2", x"3c2", x"3cf", x"3e1", x"3ef", x"3f1", x"3e9", x"3d9", x"3c3", x"3ae", x"394", x"37f", x"360", 
--			x"34e", x"343", x"331", x"326", x"319", x"313", x"30c", x"30c", x"308", x"2f4", x"2e6", x"2d9", x"2de", x"300", x"32e", x"354", 
--			x"374", x"385", x"390", x"397", x"398", x"3a5", x"3b6", x"3da", x"3f6", x"401", x"40a", x"418", x"417", x"40e", x"3ed", x"3bd", 
--			x"38b", x"361", x"33d", x"31a", x"2fd", x"2ef", x"2eb", x"2f6", x"2f7", x"2fc", x"2f7", x"2f7", x"2fc", x"2f9", x"2fe", x"303", 
--			x"310", x"315", x"31f", x"324", x"32f", x"340", x"357", x"379", x"395", x"3b2", x"3cc", x"3e0", x"3f8", x"408", x"40f", x"412", 
--			x"40f", x"40a", x"405", x"3fa", x"3e1", x"3c5", x"3a6", x"394", x"3a1", x"3c4", x"3ea", x"3ff", x"419", x"432", x"44d", x"463", 
--			x"478", x"48d", x"4a4", x"4af", x"4a6", x"494", x"473", x"454", x"43a", x"40f", x"3de", x"3b0", x"384", x"371", x"364", x"356", 
--			x"352", x"353", x"34b", x"349", x"345", x"33b", x"329", x"321", x"326", x"32f", x"33d", x"345", x"352", x"352", x"339", x"32b", 
--			x"323", x"335", x"35a", x"379", x"394", x"3b1", x"3cb", x"3d7", x"3d0", x"3c0", x"3b9", x"3c3", x"3cb", x"3e0", x"3f5", x"3f9", 
--			x"404", x"40c", x"413", x"416", x"411", x"3fd", x"3dd", x"3bb", x"39e", x"383", x"371", x"360", x"356", x"356", x"358", x"360", 
--			x"36a", x"372", x"37a", x"388", x"393", x"3a5", x"3be", x"3d0", x"3d8", x"3d2", x"3c8", x"3b2", x"395", x"385", x"37e", x"370", 
--			x"361", x"353", x"345", x"335", x"32e", x"322", x"313", x"307", x"312", x"31d", x"332", x"341", x"34c", x"353", x"357", x"35c", 
--			x"362", x"364", x"370", x"379", x"379", x"380", x"385", x"380", x"380", x"375", x"366", x"35b", x"351", x"350", x"362", x"37e", 
--			x"3b0", x"3dd", x"411", x"433", x"442", x"441", x"42f", x"400", x"3c2", x"381", x"35b", x"346", x"34c", x"36a", x"398", x"3d0", 
--			x"3fc", x"41d", x"429", x"419", x"406", x"401", x"402", x"3fc", x"3f3", x"3d7", x"3b9", x"39d", x"394", x"38f", x"389", x"386", 
--			x"386", x"385", x"394", x"39c", x"3b0", x"3b5", x"3c2", x"3c8", x"3b0", x"393", x"374", x"35f", x"34b", x"338", x"325", x"31c", 
--			x"310", x"30c", x"2fb", x"2dc", x"2ca", x"2c0", x"2b9", x"2be", x"2c5", x"2ce", x"2d9", x"2dd", x"2d6", x"2c9", x"2c5", x"2c9", 
--			x"2cf", x"2d7", x"2e1", x"2f4", x"30a", x"31a", x"32e", x"33b", x"345", x"34a", x"344", x"341", x"339", x"335", x"338", x"33f", 
--			x"345", x"350", x"355", x"35c", x"366", x"36d", x"371", x"37d", x"379", x"371", x"361", x"34c", x"332", x"31d", x"313", x"30a", 
--			x"2fb", x"2f1", x"2e7", x"2e2", x"2e6", x"2f2", x"302", x"30d", x"31a", x"320", x"31c", x"313", x"310", x"315", x"312", x"315", 
--			x"312", x"313", x"30c", x"30d", x"30a", x"314", x"31f", x"32d", x"331", x"33a", x"333", x"331", x"333", x"32f", x"333", x"338", 
--			x"33a", x"33e", x"33a", x"335", x"335", x"337", x"338", x"343", x"348", x"350", x"356", x"356", x"35a", x"35d", x"360", x"35e", 
--			x"35f", x"35c", x"355", x"358", x"35f", x"362", x"36d", x"373", x"379", x"381", x"38a", x"395", x"399", x"39e", x"39e", x"397", 
--			x"390", x"389", x"385", x"383", x"381", x"381", x"384", x"388", x"387", x"38c", x"399", x"3a3", x"3b1", x"3b8", x"3bc", x"3b6", 
--			x"3b4", x"3af", x"3a9", x"3a6", x"3a2", x"396", x"397", x"390", x"392", x"38c", x"38a", x"38a", x"38c", x"390", x"392", x"38b", 
--			x"383", x"381", x"377", x"372", x"370", x"36b", x"364", x"361", x"359", x"354", x"352", x"34f", x"354", x"353", x"351", x"34f", 
--			x"34f", x"347", x"343", x"336", x"32b", x"322", x"31d", x"31e", x"320", x"326", x"32d", x"327", x"328", x"321", x"321", x"325", 
--			x"32b", x"32f", x"335", x"335", x"33c", x"33c", x"33d", x"344", x"34a", x"355", x"35b", x"369", x"371", x"381", x"397", x"3a4", 
--			x"3b9", x"3cc", x"3d9", x"3dd", x"3e1", x"3ed", x"3f1", x"3f6", x"3fb", x"402", x"405", x"406", x"40d", x"40f", x"417", x"420", 
--			x"423", x"41d", x"420", x"417", x"41a", x"416", x"414", x"413", x"40f", x"40e", x"40e", x"40f", x"412", x"41b", x"41e", x"420", 
--			x"423", x"41d", x"41e", x"41c", x"419", x"41a", x"415", x"413", x"40c", x"401", x"3fc", x"3f9", x"3f5", x"3f3", x"3f0", x"3ef", 
--			x"3e5", x"3e0", x"3dc", x"3d2", x"3d4", x"3cf", x"3d0", x"3cd", x"3c8", x"3c4", x"3c1", x"3c1", x"3bf", x"3c5", x"3c6", x"3c5", 
--			x"3c5", x"3c1", x"3c1", x"3bd", x"3be", x"3ba", x"3b4", x"3b4", x"3af", x"3a8", x"3a2", x"3a0", x"39a", x"393", x"38e", x"38e", 
--			x"38a", x"38e", x"38a", x"38d", x"388", x"383", x"37e", x"37b", x"376", x"372", x"36b", x"36c", x"36c", x"36c", x"371", x"377", 
--			x"37a", x"37a", x"37d", x"37c", x"37e", x"386", x"384", x"38b", x"385", x"387", x"388", x"384", x"385", x"381", x"384", x"383", 
--			x"381", x"38a", x"389", x"38d", x"392", x"38f", x"392", x"38f", x"391", x"394", x"39a", x"39b", x"3ad", x"3af", x"3b1", x"3ab", 
--			x"3af", x"3ac", x"3ab", x"3a9", x"3a2", x"3b0", x"3a5", x"3ae", x"3a7", x"3a6", x"3a3", x"3a5", x"3a3", x"3ad", x"3b0", x"3ae", 
--			x"3ad", x"3ac", x"3aa", x"3a5", x"3a3", x"3a4", x"39d", x"3a5", x"3a5", x"3a6", x"3a6", x"3ab", x"3a8", x"3af", x"3ac", x"3b0", 
--			x"3ad", x"3ac", x"3ab", x"3aa", x"3ad", x"3ad", x"3a4", x"3a7", x"3ae", x"3a6", x"3ad", x"3aa", x"3a5", x"39f", x"3a0", x"39f", 
--			x"3a0", x"3a8", x"3a5", x"3ac", x"3a5", x"3a9", x"3a3", x"3a3", x"3a3", x"39e", x"3a4", x"3ae", x"3a5", x"3a7", x"3a4", x"3a5", 
--			x"3a8", x"3a7", x"3a5", x"39f", x"3ab", x"3a5", x"3a1", x"3a4", x"39f", x"39a", x"3a2", x"3a4", x"3a2", x"3a0", x"3a3", x"399", 
--			x"3a2", x"3a2", x"3a3", x"3a5", x"3a0", x"3a0", x"3a4", x"39e", x"39e", x"39e", x"3a1", x"3a0", x"3a3", x"39f", x"39e", x"3a0", 
--			x"39b", x"398", x"39a", x"39e", x"39d", x"3a3", x"39d", x"39b", x"39a", x"39c", x"39a", x"393", x"39e", x"39c", x"399", x"395", 
--			x"395", x"394", x"39c", x"39e", x"39b", x"39d", x"3a0", x"3a1", x"39c", x"39e", x"39d", x"39d", x"3a1", x"39d", x"395", x"394", 
--			x"393", x"39a", x"39a", x"3a2", x"3a4", x"3a7", x"39b", x"398", x"3a2", x"39c", x"398", x"39e", x"3a2", x"399", x"399", x"3a1", 
--			x"39c", x"398", x"39f", x"39d", x"3a0", x"3a5", x"39e", x"39e", x"3a1", x"39f", x"39e", x"3a4", x"3a2", x"3a4", x"3a1", x"39e", 
--			x"39d", x"39f", x"3a0", x"3a3", x"3a5", x"39a", x"39c", x"39f", x"399", x"39e", x"3a0", x"3a6", x"39f", x"39f", x"3a2", x"39d", 
--			x"3a1", x"3a4", x"39e", x"396", x"39f", x"39b", x"3a2", x"3a2", x"3a6", x"3a7", x"3a6", x"3a4", x"3a5", x"3a4", x"3a3", x"3a1", 
--			x"399", x"3a1", x"39c", x"39c", x"3a2", x"3a3", x"39d", x"39e", x"39e", x"39e", x"3a6", x"39e", x"3a2", x"3a7", x"3a8", x"3a5", 
--			x"39e", x"3a3", x"3a1", x"3a1", x"3a2", x"3a5", x"3a1", x"3a5", x"3a1", x"3a3", x"3a3", x"3a3", x"3aa", x"3aa", x"3aa", x"3a5", 
--			x"39f", x"3a1", x"3a6", x"3a5", x"3a6", x"3a4", x"3a6", x"39f", x"39a", x"39b", x"3a1", x"3ad", x"3a5", x"3a9", x"3a5", x"3a0", 
--			x"3a0", x"3a6", x"3a7", x"3a1", x"3ac", x"3a1", x"3a1", x"3a2", x"3a4", x"3aa", x"3a8", x"3a5", x"3a1", x"3a8", x"3a8", x"3a2", 
--			x"3aa", x"3a3", x"3a3", x"3a5", x"3aa", x"3a7", x"3a9", x"3a1", x"3a0", x"39f", x"3a1", x"3a4", x"3a9", x"3a5", x"3a3", x"3a5", 
--			x"3a4", x"39f", x"3a2", x"3ac", x"3a9", x"3ad", x"3a3", x"3a9", x"3a2", x"3a3", x"39d", x"3a8", x"3a1", x"3a2", x"3a9", x"3a3", 
--			x"3a6", x"3a5", x"3a5", x"3ae", x"3aa", x"3a3", x"3ac", x"3a7", x"3a3", x"3a0", x"3a6", x"3a3", x"3a3", x"3a1", x"3a4", x"3a3", 
--			x"3a1", x"39e", x"3a8", x"3ab", x"3a5", x"3a2", x"3aa", x"3a2", x"3a0", x"3a3", x"39d", x"39a", x"3a2", x"3a8", x"3a3", x"3a4", 
--			x"3a5", x"3a4", x"3a6", x"3ab", x"3ab", x"3a7", x"3a1", x"3aa", x"3a3", x"3a2", x"3a1", x"39e", x"39d", x"3a5", x"39e", x"39d", 
--			x"3a5", x"39d", x"3a4", x"3a7", x"3aa", x"3a9", x"3aa", x"3ad", x"3a7", x"3ab", x"39e", x"39b", x"39b", x"3a1", x"3a1", x"39f", 
--			x"3a2", x"39e", x"3a1", x"3a6", x"3ab", x"3a7", x"3a6", x"3aa", x"3a6", x"3a3", x"3a2", x"3a0", x"39f", x"3a7", x"39f", x"39f", 
--			x"39f", x"39a", x"39e", x"3a0", x"3a3", x"39e", x"3a4", x"3a5", x"3a6", x"3a5", x"3a4", x"3a3", x"3a2", x"39d", x"39e", x"39c", 
--			x"3a2", x"3a1", x"3a8", x"3a8", x"3af", x"3a3", x"3a2", x"3a5", x"3a4", x"3a8", x"3a7", x"3aa", x"3a1", x"3aa", x"3a1", x"39e", 
--			x"39e", x"39d", x"3a4", x"3a6", x"3a9", x"3a8", x"3ae", x"3aa", x"3a9", x"3ad", x"3ac", x"3ab", x"3b2", x"3ac", x"3a9", x"3a4", 
--			x"3a6", x"3a4", x"3ad", x"3a1", x"3aa", x"3a7", x"3a3", x"3a5", x"3a7", x"3ad", x"3aa", x"3ab", x"3b2", x"3b2", x"3a9", x"3a2", 
--			x"3a8", x"3a3", x"3a7", x"3a8", x"3b0", x"3af", x"3a8", x"3a6", x"3a3", x"3a1", x"3a2", x"3a9", x"3a7", x"3a6", x"3a5", x"3ac", 
--			x"3a9", x"3a8", x"3a5", x"3a5", x"3a5", x"3a2", x"3a2", x"3a5", x"3a7", x"3a9", x"3a9", x"3ac", x"3a8", x"3a9", x"3ad", x"3ac", 
--			x"3ac", x"3a9", x"3a8", x"3a2", x"3a9", x"3a5", x"3a7", x"3aa", x"3a9", x"3aa", x"3b2", x"3a8", x"3b3", x"3b3", x"3b1", x"3ae", 
--			x"3a8", x"3a8", x"3ad", x"3ad", x"3a3", x"3a9", x"3a6", x"3aa", x"3a3", x"3a5", x"3ac", x"3b3", x"3b2", x"3b1", x"3b0", x"3a7", 
--			x"3a5", x"3ac", x"3ac", x"3aa", x"3a7", x"3a9", x"3a9", x"3a8", x"3b2", x"3a4", x"3b0", x"3ad", x"3ad", x"3ab", x"3ac", x"3ad", 
--			x"3ab", x"3ab", x"3ae", x"3a9", x"3ad", x"3af", x"3a8", x"3ab", x"3aa", x"3aa", x"3a7", x"3a5", x"3ae", x"3af", x"3ae", x"3af", 
--			x"3b3", x"3a9", x"3af", x"3aa", x"3b2", x"3ab", x"3ab", x"3aa", x"3a6", x"3a5", x"3a7", x"3aa", x"3ac", x"3a6", x"3ab", x"3ac", 
--			x"3a8", x"3ad", x"3ad", x"3ac", x"3ae", x"3a5", x"3a6", x"3aa", x"3a5", x"3a9", x"3a1", x"3a3", x"3a2", x"3ac", x"3ae", x"3ae", 
--			x"3b0", x"3b0", x"3b2", x"3a8", x"3ac", x"3aa", x"39e", x"3a9", x"3a9", x"3a6", x"3a8", x"3ac", x"3b0", x"3b3", x"3a9", x"3ad", 
--			x"3a9", x"3a5", x"3ac", x"3ad", x"3ae", x"3ae", x"3ac", x"3a6", x"3a9", x"3a8", x"3a0", x"3ae", x"3a5", x"3a7", x"3aa", x"3aa", 
--			x"3ac", x"3b2", x"3ad", x"3ac", x"3b2", x"3ad", x"3ae", x"3a9", x"3a9", x"3a5", x"3ac", x"3a9", x"3a9", x"3aa", x"3a3", x"3a5", 
--			x"3a7", x"3aa", x"3a9", x"3ab", x"3b3", x"3ad", x"3ad", x"3b1", x"3a6", x"3a4", x"3a5", x"3aa", x"3aa", x"3ad", x"3ac", x"3ad", 
--			x"3aa", x"3a8", x"3b4", x"3b3", x"3b3", x"3ad", x"3ad", x"3b1", x"3ae", x"3b1", x"3ad", x"3ab", x"3a5", x"3ac", x"3ab", x"3a9", 
--			x"3af", x"3a8", x"3b0", x"3ae", x"3b0", x"3b2", x"3ae", x"3b1", x"3ad", x"3a6", x"3a9", x"3ae", x"3a8", x"3aa", x"3aa", x"3a9", 
--			x"3a6", x"3ab", x"3ab", x"3ad", x"3af", x"3a9", x"3b1", x"3b2", x"3b0", x"3ad", x"3ad", x"3a3", x"3aa", x"3a3", x"3a8", x"3a5", 
--			x"3a4", x"3a8", x"3a4", x"3aa", x"3af", x"3a8", x"3ae", x"3a3", x"3ab", x"3a7", x"3a6", x"3a4", x"3ad", x"3a5", x"3a3", x"3a5", 
--			x"39d", x"39e", x"3a3", x"3a0", x"3ae", x"3a9", x"3ad", x"3ac", x"3a5", x"3ab", x"3a3", x"3ae", x"3a6", x"3a5", x"3a5", x"39e", 
--			x"3a2", x"3a6", x"3a5", x"3a5", x"3a3", x"3a4", x"3a6", x"39e", x"3a7", x"3a6", x"3ab", x"3a6", x"3a6", x"3a5", x"3a3", x"3a3", 
--			x"3a1", x"3a0", x"3a4", x"3a4", x"3a8", x"3a1", x"3a3", x"3a4", x"3ac", x"3ab", x"3a9", x"3ad", x"3a7", x"3a6", x"3ac", x"3a6", 
--			x"3aa", x"3a5", x"3a5", x"3ab", x"3a5", x"3a5", x"3a1", x"3a2", x"3a6", x"3a6", x"3a5", x"3a7", x"3a9", x"3ab", x"3a8", x"3a2", 
--			x"3a1", x"3a2", x"3a3", x"3aa", x"3a9", x"3a4", x"3a8", x"3a7", x"3a1", x"3a8", x"3a5", x"3a4", x"3ad", x"3a9", x"3ad", x"3ac", 
--			x"3a6", x"3a2", x"3a9", x"3a4", x"3a3", x"3a1", x"3ac", x"3a3", x"39d", x"3a3", x"3a9", x"3ae", x"3b0", x"3b3", x"3a4", x"3ab", 
--			x"3a6", x"3a7", x"3a4", x"3a5", x"3a9", x"3a7", x"3ac", x"3a8", x"3a1", x"3a7", x"3a5", x"3aa", x"3a9", x"3aa", x"3ad", x"3aa", 
--			x"3b2", x"3a7", x"3a6", x"3a8", x"3a7", x"3a6", x"3a8", x"3ac", x"3a9", x"3ad", x"3b0", x"3a9", x"3ad", x"3a6", x"3a8", x"3a2", 
--			x"3a6", x"3b2", x"3b1", x"3b2", x"3ac", x"3ab", x"3aa", x"3a8", x"3a1", x"3a7", x"3ac", x"3ac", x"3ac", x"3af", x"3ab", x"3a9", 
--			x"3a9", x"3aa", x"3af", x"3b0", x"3af", x"3a9", x"3a4", x"3b0", x"3a6", x"3a0", x"3ad", x"3a8", x"3a5", x"3a2", x"3a5", x"3a9", 
--			x"3a3", x"3ac", x"3ab", x"3a6", x"3a8", x"3aa", x"3a9", x"3a6", x"3a4", x"3a4", x"3aa", x"3a1", x"3a3", x"3a3", x"3a8", x"3a7", 
--			x"3aa", x"3a3", x"3ab", x"3a4", x"3a5", x"3a5", x"3aa", x"3a9", x"3a5", x"3a6", x"3a9", x"3a6", x"3a3", x"3a7", x"3ae", x"3a6", 
--			x"3a8", x"3ad", x"3a4", x"3ae", x"3ab", x"3a6", x"3ae", x"3a9", x"3ad", x"3ac", x"3a9", x"3a7", x"3ac", x"3aa", x"3ac", x"3ae", 
--			x"3ac", x"3ab", x"3ae", x"3ad", x"3ab", x"3ad", x"3ad", x"3ac", x"3ac", x"3b2", x"3b1", x"3a9", x"3b4", x"3ae", x"3a7", x"3aa", 
--			x"3b0", x"3ae", x"3a8", x"3ab", x"3b0", x"3ab", x"3ae", x"3ab", x"3a5", x"3ae", x"3b1", x"3ac", x"3ad", x"3a9", x"3a8", x"3a1", 
--			x"3aa", x"3ae", x"3a8", x"3b1", x"3ad", x"3ad", x"3ad", x"3b1", x"3b2", x"3ab", x"3aa", x"3a5", x"3a5", x"3a8", x"3a8", x"3ad", 
--			x"3a2", x"3ab", x"3a5", x"3aa", x"3a8", x"3a9", x"3aa", x"3a5", x"3a9", x"3ae", x"3ac", x"3b0", x"3a9", x"3aa", x"3a5", x"3a6", 
--			x"3a0", x"3a8", x"3a6", x"3a5", x"3aa", x"3a6", x"3ac", x"3a9", x"3ac", x"3a8", x"3ab", x"3a5", x"3a7", x"3aa", x"3ac", x"3a6", 
--			x"3b0", x"3a9", x"3ad", x"3a4", x"3aa", x"3a9", x"3a8", x"3a9", x"3ae", x"3a8", x"3aa", x"3ab", x"3ab", x"3a6", x"3a6", x"3a9", 
--			x"3aa", x"3a0", x"3ab", x"3a3", x"3a9", x"3a4", x"3a9", x"3aa", x"3a9", x"3a8", x"3a8", x"3a4", x"3a6", x"3ab", x"3a2", x"3a8", 
--			x"3a1", x"3ab", x"3a9", x"3a8", x"3a4", x"3ae", x"3a3", x"3a5", x"3ab", x"3a5", x"3a1", x"3a9", x"3ab", x"3aa", x"3a1", x"3ac", 
--			x"3ad", x"3aa", x"3a1", x"3ab", x"3aa", x"3ac", x"3ac", x"3a9", x"3ae", x"3ae", x"3a6", x"3ae", x"3ad", x"3a7", x"3ad", x"3ae", 
--			x"3ac", x"3af", x"3a7", x"3ae", x"3aa", x"3ab", x"3a6", x"3ab", x"3a9", x"3ad", x"3ad", x"3a9", x"3aa", x"3ad", x"3ac", x"3af",
--			x"3b6", x"3ad", x"3a8", x"3ad", x"3b0", x"3ab", x"3a7", x"3aa", x"3a9", x"3ad", x"3b1", x"3a6", x"3ab", x"3ab", x"3a5", x"3a9", 
--			x"3ac", x"3af", x"3aa", x"3ae", x"3a8", x"3ad", x"3a9", x"3a8", x"3ab", x"3a5", x"3ad", x"3a8", x"3a9", x"3a8", x"3b3", x"3a7", 
--			x"3a6", x"3ae", x"3ab", x"3b1", x"3aa", x"3a6", x"3a6", x"3ad", x"3ab", x"3a6", x"3ad", x"3a9", x"3ae", x"3af", x"3ae", x"3aa", 
--			x"3ab", x"3ad", x"3af", x"3ac", x"3b0", x"3af", x"3af", x"3ad", x"3b2", x"3b6", x"3b1", x"3b4", x"3b5", x"3b0", x"3b1", x"3ad", 
--			x"3b2", x"3aa", x"3a7", x"3b0", x"3af", x"3af", x"3ad", x"3b4", x"3ad", x"3ac", x"3b2", x"3ac", x"3ba", x"3b3", x"3b2", x"3ba", 
--			x"3b6", x"3b5", x"3ad", x"3af", x"3b4", x"3b3", x"3b2", x"3b3", x"3b2", x"3af", x"3a9", x"3b4", x"3b2", x"3ad", x"3b2", x"3ab", 
--			x"3b0", x"3aa", x"3b2", x"3b0", x"3b2", x"3ad", x"3ad", x"3ac", x"3b0", x"3aa", x"3ac", x"3a6", x"3af", x"3ae", x"3ab", x"3ad", 
--			x"3ab", x"3af", x"3a3", x"3aa", x"3ab", x"3a7", x"3a6", x"3a8", x"3ad", x"3af", x"3ac", x"3b1", x"3b1", x"3ae", x"3af", x"3a9", 
--			x"3ad", x"3a9", x"3ad", x"3ad", x"3b0", x"3a9", x"3ac", x"3ad", x"3a9", x"3ac", x"3ac", x"3b6", x"3af", x"3b0", x"3ad", x"3aa", 
--			x"3b2", x"3ad", x"3a8", x"3a9", x"3ac", x"3aa", x"3ad", x"3ad", x"3ae", x"3a5", x"3a5", x"3a7", x"3a4", x"3ad", x"3a7", x"3a4", 
--			x"3aa", x"3a9", x"3aa", x"3a9", x"3a8", x"3aa", x"3a2", x"3a5", x"3a9", x"3a7", x"3a3", x"3a7", x"3a6", x"3ab", x"3a1", x"3a7", 
--			x"3aa", x"3a7", x"3a5", x"3a2", x"3ab", x"3a9", x"3aa", x"3ac", x"3aa", x"3a3", x"3a8", x"3aa", x"3ae", x"3ac", x"3a8", x"3af", 
--			x"3a5", x"3a7", x"3a9", x"3ad", x"3ad", x"3ab", x"3ab", x"39f", x"3a7", x"3ad", x"3ad", x"3a9", x"3a1", x"3ae", x"3ab", x"3a6", 
--			x"3aa", x"3b2", x"3b1", x"3af", x"3b4", x"3b0", x"3af", x"3af", x"3af", x"3ad", x"3ac", x"3b0", x"3ae", x"3ad", x"3ac", x"3b0", 
--			x"3a9", x"3ab", x"3af", x"3ae", x"3ab", x"3ab", x"3af", x"3a1", x"3a6", x"3a6", x"3a7", x"3a4", x"3a3", x"3a4", x"3b0", x"3ab", 
--			x"3a5", x"3a4", x"3a4", x"3aa", x"3a1", x"3a6", x"3a6", x"3a6", x"3a4", x"3a6", x"3a1", x"3aa", x"3a4", x"3a9", x"3a7", x"3a5",
--			x"3a4", x"3a9", x"3a4", x"3b0", x"3a9", x"39d", x"3a9", x"3a7", x"3a7", x"3a7", x"3a9", x"3a1", x"3aa", x"3ad", x"3a5", x"3a3", 
--			x"3a6", x"3ab", x"3a7", x"3a8", x"3a6", x"3a2", x"3a8", x"3b0", x"3b0", x"3ab", x"3a6", x"3a3", x"3aa", x"3b1", x"3ac", x"3a8", 
--			x"3ac", x"3b4", x"3ae", x"3ad", x"3a7", x"3ac", x"3ac", x"3aa", x"3ac", x"3ad", x"3a8", x"3ad", x"3b0", x"3ad", x"3a9", x"3a9", 
--			x"3b3", x"3ab", x"3a6", x"3ae", x"3aa", x"3ae", x"3af", x"3b0", x"3b2", x"3ab", x"3a8", x"3a5", x"3ad", x"3ac", x"3a7", x"3a3", 
--			x"3a8", x"3a6", x"3ae", x"3a3", x"3a1", x"3a0", x"3ad", x"3ae", x"3aa", x"3a3", x"3a7", x"3a2", x"3a9", x"3a4", x"399", x"39f", 
--			x"3a7", x"3a9", x"3a5", x"3a3", x"3a8", x"3ad", x"3ae", x"3aa", x"3a6", x"39e", x"3a6", x"3ae", x"3ac", x"3aa", x"3a1", x"3aa", 
--			x"3a8", x"3a6", x"3a4", x"3a0", x"3a7", x"3a4", x"3ac", x"3a4", x"39e", x"39a", x"39a", x"39a", x"39f", x"39b", x"3a2", x"3ab", 
--			x"3a4", x"3a8", x"3a2", x"39b", x"399", x"395", x"399", x"39e", x"39f", x"3ad", x"3a4", x"3a8", x"3a1", x"3a9", x"3a7", x"3a3", 
--			x"3a8", x"3b4", x"3b8", x"3b7", x"3ae", x"3a4", x"3a4", x"3a2", x"3a5", x"3a9", x"39c", x"3a7", x"3a0", x"3aa", x"3b3", x"39a", 
--			x"39d", x"38b", x"397", x"39a", x"3a3", x"39d", x"3a3", x"39e", x"39f", x"397", x"38f", x"388", x"39a", x"396", x"39b", x"3a7", 
--			x"3a8", x"3a5", x"3a8", x"3a2", x"39d", x"39b", x"39d", x"3a1", x"3a5", x"3a2", x"3a1", x"3aa", x"3c0", x"3c8", x"3b8", x"3a0", 
--			x"3a3", x"39d", x"3a1", x"3a3", x"3a5", x"3ab", x"3b7", x"3b9", x"3b1", x"3a6", x"39e", x"39f", x"3a0", x"3ab", x"3aa", x"3aa", 
--			x"3a4", x"39f", x"39e", x"3a0", x"3a8", x"3aa", x"3b8", x"3b1", x"3af", x"3ae", x"39e", x"39b", x"39b", x"396", x"395", x"39f", 
--			x"3ab", x"3c2", x"3b9", x"3b5", x"3a6", x"3a4", x"3a2", x"3a0", x"399", x"39e", x"3b0", x"3b0", x"3a2", x"3a6", x"3b1", x"3bb", 
--			x"3bc", x"3b0", x"3b0", x"39f", x"3a6", x"3a1", x"3a4", x"39d", x"3a3", x"3a5", x"3b8", x"3b8", x"3ad", x"3a8", x"3b1", x"3bf", 
--			x"3c8", x"3bd", x"3b1", x"3ae", x"3bf", x"3af", x"3a7", x"3a7", x"3b4", x"3c6", x"3c9", x"3b5", x"3ab", x"3a0", x"3a0", x"3a3",
--			x"398", x"399", x"39c", x"3a9", x"3b2", x"3aa", x"39d", x"393", x"39a", x"3ab", x"3a9", x"3ad", x"3ba", x"3ba", x"3c1", x"3cf", 
--			x"3c0", x"3b9", x"3b3", x"3b1", x"3b5", x"3b1", x"3af", x"3b1", x"3c4", x"3cb", x"3bd", x"3b1", x"3af", x"3aa", x"3a8", x"3b3", 
--			x"3b1", x"3bf", x"3c7", x"3c5", x"3d6", x"3c6", x"3bb", x"3a2", x"393", x"397", x"3a7", x"3b2", x"3bd", x"3cc", x"3df", x"3e2", 
--			x"3d8", x"3b3", x"383", x"37f", x"385", x"3a4", x"3c1", x"3b4", x"3ae", x"3b0", x"3aa", x"3ab", x"3a6", x"393", x"399", x"3b7", 
--			x"3c9", x"3bf", x"3a4", x"39d", x"395", x"3a3", x"3a9", x"3b3", x"3ac", x"3bd", x"3cb", x"3ca", x"3bd", x"3b5", x"3ac", x"3a8", 
--			x"39f", x"39c", x"3aa", x"3af", x"3c0", x"3c0", x"3c1", x"3c2", x"3b9", x"3ac", x"39e", x"39f", x"398", x"3a4", x"3a0", x"39f", 
--			x"396", x"3a8", x"3b5", x"3b6", x"3af", x"3a3", x"3a1", x"3ab", x"3b0", x"3ab", x"39c", x"399", x"399", x"3b0", x"3af", x"3a4", 
--			x"3a4", x"3af", x"3b5", x"3c1", x"3b4", x"3a6", x"39e", x"3b3", x"3b9", x"3b7", x"3b1", x"3ac", x"3ac", x"3b6", x"3b3", x"3ac"
--			);

		constant DATA_ROM : ROM := (
			x"3a9", x"3af", x"3aa", x"3a7", x"3a7", x"3aa", x"3aa", x"3b0", x"3a4", x"3a8", x"3a3", x"3a0", x"3a1", x"39d", x"3a3", x"3a3", 
			x"3ac", x"3a8", x"3a5", x"3a5", x"3a1", x"3a8", x"3a3", x"3a0", x"398", x"3a5", x"3a3", x"3a6", x"3ae", x"3aa", x"3ae", x"3ac", 
			x"3a5", x"3a4", x"3a1", x"3a7", x"3aa", x"3a3", x"3a9", x"3aa", x"3a2", x"3a4", x"3a5", x"39f", x"3a6", x"3aa", x"3ac", x"3ac", 
			x"3a8", x"3ac", x"3ac", x"3a6", x"3ab", x"3aa", x"3a9", x"3a9", x"3ac", x"3ac", x"3a7", x"3a5", x"3a7", x"3a7", x"3ab", x"3a5", 
			x"3a5", x"39f", x"39f", x"3a3", x"39f", x"39c", x"3a4", x"3a0", x"3ae", x"3aa", x"3b2", x"3af", x"3aa", x"3a3", x"3a9", x"3a0", 
			x"3a1", x"3aa", x"3ac", x"3ad", x"3a7", x"3af", x"3a5", x"3ab", x"3a8", x"3a7", x"3a2", x"3a0", x"3a3", x"3a7", x"3ab", x"3a3", 
			x"3ab", x"3a6", x"3a5", x"3aa", x"3ad", x"3a5", x"3ab", x"3b3", x"3aa", x"3ae", x"3aa", x"3aa", x"3a5", x"3a1", x"3a6", x"3a5", 
			x"3a4", x"3b0", x"3a2", x"3a2", x"3a9", x"3a5", x"3a2", x"3a3", x"3a3", x"3a4", x"39f", x"3a1", x"3a3", x"3a0", x"3a6", x"3a1", 
			x"3a6", x"3ac", x"3ac", x"3ac", x"3a8", x"3a8", x"3a8", x"3a5", x"3b1", x"3af", x"3ab", x"3aa", x"3b2", x"3a5", x"3ab", x"3b3", 
			x"3a9", x"396", x"3c1", x"3bb", x"3a8", x"3a2", x"3a8", x"38f", x"3b4", x"3cc", x"38a", x"3b1", x"3ae", x"38a", x"3b9", x"3bb", 
			x"3a0", x"3af", x"3a7", x"39b", x"3b1", x"3c3", x"3ab", x"3a9", x"3a8", x"395", x"3b5", x"3bd", x"3a3", x"3af", x"3af", x"3a1", 
			x"3ab", x"3bc", x"3a7", x"3a9", x"3af", x"39c", x"39e", x"3b6", x"3a4", x"3a6", x"3a4", x"39c", x"39d", x"3a8", x"3a1", x"39c", 
			x"3a8", x"3a0", x"3a1", x"3ad", x"39f", x"39f", x"3a9", x"39e", x"39f", x"3ad", x"3a3", x"395", x"3a1", x"399", x"395", x"3ab", 
			x"3a7", x"3a6", x"39b", x"39d", x"39d", x"39d", x"39f", x"3a6", x"3ac", x"3a8", x"39f", x"3a8", x"3ab", x"39f", x"3a3", x"3a0", 
			x"39d", x"39f", x"3a5", x"39f", x"3ac", x"3a3", x"39d", x"3ab", x"3a9", x"3a3", x"3a0", x"3a8", x"3a5", x"3a8", x"3a8", x"3a6", 
			x"3a3", x"3a8", x"3ab", x"3a7", x"3a9", x"3aa", x"3a3", x"3a5", x"3a5", x"3a9", x"3ad", x"3a9", x"3ae", x"3a9", x"3a5", x"3ae", 
			x"3a7", x"3af", x"3aa", x"3ad", x"3ab", x"3a0", x"3a2", x"3a5", x"3a1", x"39e", x"3a3", x"3a9", x"3a5", x"3a3", x"39d", x"3a5", 
			x"39d", x"3a2", x"3a0", x"397", x"399", x"3a4", x"3ac", x"3ac", x"3a3", x"398", x"3a3", x"3a9", x"39c", x"3a0", x"3a5", x"39d", 
			x"3a2", x"3a2", x"39f", x"3a9", x"3a6", x"3a5", x"39f", x"3a2", x"3a9", x"3ac", x"3a5", x"3a2", x"39a", x"3ad", x"3a7", x"3a5", 
			x"3a2", x"39d", x"3a4", x"3a7", x"3a4", x"3aa", x"3a3", x"3a5", x"3ad", x"3a1", x"3a7", x"3b9", x"3b7", x"3bb", x"3b3", x"3b7", 
			x"3b6", x"3b7", x"3ba", x"3b6", x"3b2", x"3b4", x"3b5", x"3b5", x"3b8", x"3b8", x"3b3", x"3ba", x"3b1", x"3b5", x"3b9", x"3b5", 
			x"3b2", x"3b3", x"3b5", x"3b2", x"3b1", x"3b3", x"3b7", x"3ae", x"3b3", x"3b0", x"3b2", x"3ac", x"3ab", x"3b1", x"3af", x"3af", 
			x"3ad", x"3b1", x"3ad", x"3a5", x"3ad", x"3b1", x"3ac", x"3a4", x"3a0", x"3a2", x"39e", x"3a0", x"3aa", x"3a4", x"3a3", x"39f", 
			x"39b", x"3a5", x"3a4", x"3a5", x"3ad", x"3a8", x"3a8", x"3a8", x"3a4", x"3a9", x"3a8", x"3a6", x"3a0", x"39f", x"39f", x"3a4", 
			x"3a5", x"3ad", x"3ab", x"39f", x"3ab", x"3a4", x"3b2", x"3b2", x"3ac", x"3aa", x"3a9", x"3af", x"3ae", x"3a8", x"3a5", x"3a5", 
			x"3a5", x"3ac", x"3a0", x"3a8", x"3a5", x"3a6", x"3a8", x"3a4", x"39f", x"39d", x"3a8", x"3a2", x"3a4", x"3a6", x"3aa", x"3aa", 
			x"3ab", x"39b", x"39f", x"3a4", x"3a7", x"39b", x"3a3", x"39d", x"39f", x"3a3", x"3a7", x"3a7", x"39c", x"3a9", x"3a1", x"3a6", 
			x"3a8", x"3a4", x"3a8", x"3a6", x"3a0", x"3a5", x"3a3", x"3a5", x"3a9", x"39d", x"39a", x"3a3", x"3a0", x"3a2", x"3a3", x"3ab", 
			x"3a7", x"39f", x"3ab", x"3a7", x"39f", x"3ab", x"3a7", x"39f", x"3a8", x"3b3", x"3a6", x"3a2", x"3b0", x"3a9", x"3a5", x"3ae", 
			x"3ab", x"3a8", x"3a4", x"3b1", x"3ad", x"39f", x"3a8", x"3a0", x"3aa", x"3b2", x"3aa", x"39d", x"3ad", x"3b3", x"3a9", x"3a9", 
			x"3ac", x"3a9", x"3b3", x"3a3", x"3a7", x"3a8", x"3ad", x"3a7", x"3a6", x"3ad", x"3ac", x"3a9", x"3b6", x"3b2", x"3b6", x"3b6", 
			x"3b1", x"3a6", x"3b2", x"3ac", x"3a8", x"3a9", x"3a7", x"3a4", x"3ac", x"3ab", x"3a7", x"3a6", x"39d", x"3a5", x"3a8", x"3a8", 
			x"3a6", x"3a4", x"39f", x"3a8", x"3a8", x"3a5", x"3a2", x"3a1", x"39e", x"3ab", x"3ab", x"39e", x"3ac", x"3a7", x"3a1", x"3a8", 
			x"3af", x"3a6", x"3b1", x"3a3", x"3ad", x"3a5", x"3a7", x"3a0", x"3a8", x"39a", x"39b", x"39e", x"3a2", x"3a2", x"3a6", x"3a4", 
			x"3a6", x"3a5", x"39c", x"39d", x"3a6", x"3a6", x"3a2", x"3a6", x"3a5", x"39f", x"397", x"39f", x"3a6", x"3a4", x"3ab", x"3a7", 
			x"3a6", x"3ab", x"3a7", x"3a3", x"39f", x"39b", x"39b", x"3a7", x"39b", x"3a7", x"3ab", x"3aa", x"3a6", x"3a2", x"3aa", x"3a4", 
			x"3a1", x"398", x"39f", x"3a2", x"3a6", x"3a4", x"3a6", x"3a4", x"3a6", x"3a2", x"3a4", x"3a4", x"3a6", x"3a3", x"3a5", x"3a5", 
			x"3a4", x"3a8", x"39f", x"3ab", x"39c", x"3a8", x"3ad", x"3a7", x"3a9", x"3ab", x"3a4", x"3af", x"3a7", x"3a3", x"3a7", x"3a1", 
			x"3ac", x"3a9", x"3b2", x"3ac", x"3a4", x"3aa", x"3af", x"3b1", x"3a2", x"3a1", x"3a0", x"3a8", x"3aa", x"3b4", x"3a0", x"3a8", 
			x"3b4", x"3ab", x"3a8", x"3ab", x"3a7", x"3af", x"3ac", x"3af", x"3ae", x"3a9", x"3b6", x"3af", x"3ac", x"3a5", x"3a3", x"3a5", 
			x"3a3", x"3a0", x"3a3", x"3aa", x"3aa", x"3a9", x"3a6", x"3ae", x"3ae", x"3aa", x"3a7", x"3a1", x"3a4", x"3a9", x"3ac", x"3ae", 
			x"3b0", x"3b2", x"3ad", x"3b4", x"3a9", x"3b8", x"3b8", x"3c6", x"46e", x"534", x"477", x"4ab", x"386", x"340", x"368", x"391", 
			x"40e", x"432", x"41a", x"3a5", x"35f", x"38b", x"38b", x"3d3", x"411", x"3aa", x"386", x"35a", x"353", x"36c", x"3aa", x"3b0", 
			x"39e", x"38a", x"372", x"36e", x"3a6", x"405", x"47c", x"44a", x"41c", x"38a", x"339", x"33a", x"34c", x"385", x"3b6", x"3c1", 
			x"3b7", x"3a0", x"3bf", x"3cb", x"3ef", x"449", x"413", x"3a3", x"36f", x"32e", x"2f0", x"33c", x"354", x"36e", x"3a5", x"3ab", 
			x"393", x"39b", x"3ab", x"38f", x"381", x"385", x"358", x"35c", x"374", x"363", x"387", x"3a9", x"3aa", x"3ae", x"3be", x"3b6", 
			x"3be", x"3cc", x"3b6", x"39f", x"38a", x"37d", x"379", x"37f", x"38b", x"399", x"3a3", x"3af", x"3bd", x"3c3", x"3dc", x"3d9", 
			x"3f6", x"40b", x"41d", x"420", x"415", x"407", x"3d7", x"3bd", x"3c3", x"3c9", x"3dc", x"400", x"3ed", x"3de", x"3d0", x"3b8", 
			x"39d", x"38d", x"370", x"35c", x"351", x"342", x"33c", x"340", x"33c", x"32e", x"320", x"315", x"308", x"30e", x"315", x"2df", 
			x"2b1", x"284", x"2bc", x"428", x"49f", x"583", x"594", x"457", x"3f5", x"309", x"304", x"2fe", x"373", x"367", x"35b", x"36f", 
			x"36b", x"3c4", x"471", x"4c6", x"4ab", x"47d", x"3bf", x"35d", x"307", x"329", x"32f", x"37b", x"38f", x"3ad", x"441", x"50b", 
			x"522", x"54d", x"4b7", x"3e7", x"349", x"305", x"30b", x"364", x"3f5", x"41e", x"42e", x"41c", x"3d5", x"3d2", x"3d2", x"3c0", 
			x"397", x"361", x"32c", x"2ff", x"2fe", x"2f9", x"2f6", x"2d9", x"2b9", x"2b2", x"2ce", x"346", x"399", x"466", x"50f", x"4b1", 
			x"4c4", x"409", x"370", x"339", x"309", x"322", x"333", x"366", x"352", x"381", x"3cb", x"41d", x"461", x"4a9", x"46f", x"412", 
			x"3b4", x"33c", x"30c", x"30b", x"32b", x"34e", x"392", x"3c0", x"3f4", x"42d", x"47b", x"48b", x"4b7", x"49e", x"406", x"3b3", 
			x"353", x"313", x"357", x"38b", x"3e1", x"438", x"458", x"446", x"435", x"429", x"3e2", x"3c1", x"396", x"34e", x"339", x"325", 
			x"31e", x"329", x"334", x"327", x"311", x"30b", x"306", x"316", x"355", x"361", x"369", x"3a8", x"3fe", x"431", x"473", x"47e", 
			x"3f8", x"3b5", x"347", x"303", x"312", x"349", x"36c", x"3a2", x"3d3", x"3c6", x"3f3", x"41e", x"42f", x"424", x"40e", x"3a6", 
			x"34f", x"324", x"30f", x"32b", x"37e", x"3b4", x"3db", x"3f9", x"402", x"3fd", x"431", x"493", x"44f", x"44c", x"3ed", x"362", 
			x"35e", x"361", x"395", x"406", x"455", x"448", x"43b", x"418", x"3c4", x"3bc", x"3b2", x"389", x"387", x"371", x"341", x"336", 
			x"33d", x"326", x"32b", x"324", x"305", x"301", x"30e", x"301", x"326", x"342", x"352", x"390", x"434", x"461", x"494", x"4a4", 
			x"3e2", x"384", x"326", x"2da", x"302", x"34c", x"378", x"3a4", x"3d4", x"3e4", x"3fb", x"440", x"449", x"429", x"409", x"38f", 
			x"32e", x"30e", x"302", x"329", x"385", x"3c8", x"3ef", x"410", x"428", x"419", x"460", x"4a0", x"457", x"478", x"3e0", x"35b", 
			x"34a", x"31b", x"372", x"3e7", x"451", x"467", x"465", x"436", x"3c0", x"3ac", x"382", x"365", x"377", x"35d", x"343", x"344", 
			x"32d", x"321", x"32c", x"325", x"31f", x"312", x"31a", x"306", x"30a", x"335", x"358", x"3d7", x"459", x"482", x"4a1", x"44f", 
			x"3c1", x"354", x"30e", x"2fe", x"332", x"377", x"399", x"3bc", x"3d3", x"3d5", x"3fc", x"44d", x"457", x"43f", x"3f5", x"361", 
			x"315", x"2e7", x"307", x"360", x"3c3", x"411", x"422", x"42b", x"426", x"456", x"481", x"47d", x"465", x"3d6", x"36e", x"323", 
			x"319", x"381", x"3fd", x"467", x"494", x"45f", x"3f6", x"39e", x"36d", x"370", x"38d", x"3a2", x"393", x"373", x"343", x"316", 
			x"313", x"31b", x"329", x"32d", x"319", x"309", x"2f2", x"2ef", x"2f4", x"31e", x"3ab", x"473", x"49a", x"50f", x"480", x"3d8", 
			x"365", x"2d9", x"2cc", x"320", x"359", x"3a5", x"3ce", x"3cb", x"3c5", x"3df", x"41f", x"423", x"440", x"40b", x"394", x"34d", 
			x"308", x"300", x"341", x"38f", x"3dd", x"40b", x"421", x"40c", x"40e", x"440", x"46c", x"452", x"44b", x"3d8", x"363", x"34f", 
			x"33d", x"38e", x"415", x"458", x"473", x"456", x"3f4", x"3ad", x"398", x"382", x"396", x"3a8", x"395", x"375", x"355", x"333", 
			x"338", x"346", x"34b", x"345", x"329", x"30e", x"2ea", x"2e0", x"2e3", x"2de", x"2f5", x"350", x"414", x"47e", x"4f9", x"4f5", 
			x"438", x"3b9", x"30b", x"2a3", x"2e3", x"31e", x"381", x"3df", x"3e2", x"3de", x"3ca", x"3e5", x"404", x"423", x"439", x"3e8", 
			x"396", x"33f", x"2f7", x"30b", x"34c", x"3a1", x"3fe", x"431", x"431", x"41e", x"41d", x"430", x"439", x"44e", x"41a", x"3cd", 
			x"38e", x"358", x"369", x"3b1", x"3ff", x"44a", x"457", x"427", x"3e2", x"3b2", x"38f", x"3a0", x"3b8", x"3b5", x"3a6", x"37c", 
			x"349", x"331", x"334", x"344", x"360", x"363", x"345", x"31c", x"2f2", x"2dd", x"2d7", x"2d4", x"2d9", x"2f2", x"39d", x"445", 
			x"4a9", x"53b", x"4ae", x"417", x"38f", x"2c3", x"2ba", x"2ff", x"342", x"3c1", x"3fb", x"3ee", x"3d2", x"3c6", x"3de", x"401", 
			x"444", x"429", x"3d9", x"38c", x"31c", x"2e7", x"31c", x"359", x"3c1", x"427", x"441", x"43f", x"431", x"42e", x"427", x"451", 
			x"436", x"3f0", x"3bb", x"35e", x"33e", x"37c", x"3b1", x"412", x"465", x"446", x"42d", x"3e0", x"39b", x"385", x"394", x"3a3", 
			x"3ac", x"3a7", x"372", x"358", x"347", x"33f", x"356", x"365", x"355", x"33c", x"31a", x"2f1", x"2d6", x"2de", x"2d9", x"2bf", 
			x"2e0", x"37c", x"421", x"4a3", x"54b", x"4c9", x"445", x"3aa", x"2c5", x"2ba", x"2e7", x"330", x"3c4", x"409", x"3fd", x"3e3", 
			x"3bc", x"3bc", x"3e2", x"42d", x"431", x"3ff", x"3bd", x"33b", x"2fd", x"317", x"33d", x"3a8", x"414", x"43a", x"440", x"42d", 
			x"402", x"410", x"427", x"427", x"41c", x"3e7", x"392", x"37b", x"37a", x"39d", x"3fb", x"439", x"447", x"430", x"3e9", x"3a2", 
			x"386", x"380", x"39a", x"3c2", x"3cb", x"3a9", x"38c", x"35d", x"345", x"349", x"34a", x"34b", x"344", x"320", x"2fb", x"2df", 
			x"2cd", x"2cd", x"2c9", x"2c0", x"341", x"41b", x"46f", x"541", x"515", x"45c", x"3f2", x"302", x"298", x"2dd", x"303", x"38f", 
			x"3fe", x"409", x"3f1", x"3cf", x"3c9", x"3ce", x"41e", x"444", x"410", x"3e1", x"36c", x"2f7", x"309", x"310", x"367", x"3e9", 
			x"422", x"43b", x"43d", x"411", x"3e4", x"3e7", x"3f0", x"410", x"431", x"429", x"3e9", x"3ab", x"377", x"361", x"397", x"3c3", 
			x"418", x"43a", x"43b", x"411", x"3de", x"3b5", x"397", x"397", x"398", x"386", x"371", x"35d", x"33d", x"343", x"34d", x"34e", 
			x"34a", x"32a", x"2f5", x"2cf", x"2bb", x"2b8", x"2bf", x"2fc", x"3bf", x"44b", x"4bf", x"539", x"497", x"431", x"3a0", x"2d2", 
			x"2dc", x"2ee", x"32b", x"3a2", x"3e0", x"3df", x"3e8", x"3ef", x"3ff", x"410", x"465", x"417", x"3e3", x"390", x"2f6", x"2da", 
			x"2fa", x"31e", x"3a7", x"411", x"42e", x"45d", x"429", x"404", x"3d7", x"3c8", x"3a5", x"39f", x"3be", x"3b6", x"3f1", x"41b", 
			x"3ff", x"40a", x"3ec", x"39f", x"3c1", x"3a4", x"3d6", x"405", x"423", x"428", x"3fc", x"3ca", x"375", x"348", x"32e", x"32c", 
			x"352", x"37b", x"37b", x"37d", x"34f", x"312", x"2e0", x"2ba", x"2ab", x"2b0", x"2d1", x"348", x"416", x"47a", x"520", x"4f2", 
			x"45f", x"3e3", x"31e", x"2b7", x"2ee", x"312", x"396", x"3ee", x"3f5", x"3ef", x"3d0", x"3be", x"3d5", x"413", x"433", x"40e", 
			x"3d9", x"35d", x"2f1", x"2e8", x"2f5", x"360", x"3e6", x"42e", x"45b", x"44a", x"405", x"3c3", x"3a3", x"38c", x"389", x"399", 
			x"383", x"377", x"374", x"3a1", x"3e6", x"458", x"4a6", x"497", x"467", x"3f3", x"36b", x"350", x"349", x"398", x"404", x"42f", 
			x"42a", x"3ee", x"386", x"343", x"335", x"351", x"37d", x"3ab", x"395", x"35a", x"318", x"2b9", x"27f", x"26b", x"284", x"2e6", 
			x"3b3", x"47d", x"4ff", x"55b", x"4d5", x"42b", x"385", x"2cf", x"2bc", x"2ef", x"340", x"3b2", x"3ee", x"3db", x"3c5", x"3af", 
			x"3c2", x"3fb", x"44e", x"44e", x"420", x"3bc", x"325", x"2d5", x"2d1", x"2fa", x"37d", x"3ff", x"44b", x"46f", x"44e", x"40e", 
			x"3d0", x"3a6", x"383", x"37e", x"373", x"35e", x"359", x"35b", x"36d", x"3a6", x"3e8", x"43f", x"479", x"476", x"470", x"417", 
			x"3d3", x"3a2", x"364", x"37f", x"386", x"3b3", x"3da", x"3ee", x"3f4", x"3e2", x"3c4", x"3a0", x"37c", x"35d", x"345", x"330", 
			x"31d", x"302", x"2f0", x"2c1", x"2a6", x"2c5", x"323", x"3f1", x"49c", x"531", x"53f", x"4b4", x"404", x"335", x"2b7", x"2ac", 
			x"2e6", x"357", x"3bc", x"3eb", x"3e6", x"3ce", x"3c5", x"3d3", x"40d", x"435", x"42e", x"3f9", x"38a", x"320", x"2ea", x"2e3", 
			x"32a", x"39d", x"403", x"44e", x"45d", x"43a", x"3fa", x"3c3", x"393", x"379", x"36d", x"358", x"34d", x"355", x"35d", x"38a", 
			x"3bd", x"3f2", x"41f", x"425", x"417", x"3f0", x"3c3", x"396", x"379", x"366", x"377", x"396", x"3b6", x"3f5", x"3f3", x"3fa", 
			x"3f6", x"3cd", x"3c5", x"3ba", x"3b6", x"3b6", x"3bc", x"3a7", x"3a3", x"396", x"386", x"385", x"393", x"393", x"3a3", x"3ab", 
			x"39a", x"399", x"384", x"361", x"341", x"301", x"2d5", x"2c6", x"2fe", x"387", x"41e", x"4bd", x"4f2", x"49f", x"42d", x"376", 
			x"307", x"2eb", x"301", x"34f", x"397", x"3bc", x"3b6", x"3aa", x"3ac", x"3cf", x"414", x"44f", x"44e", x"425", x"3ad", x"341", 
			x"2f5", x"2db", x"313", x"374", x"3d4", x"425", x"448", x"435", x"403", x"3d7", x"3ab", x"399", x"390", x"379", x"365", x"352", 
			x"33e", x"351", x"37c", x"3c2", x"408", x"437", x"43b", x"40f", x"3cc", x"389", x"360", x"34f", x"354", x"363", x"37c", x"38a", 
			x"3a0", x"3b9", x"3da", x"3fd", x"419", x"41b", x"401", x"3d1", x"395", x"36b", x"352", x"355", x"36f", x"389", x"3a1", x"3b6", 
			x"3bd", x"3cc", x"3d7", x"3eb", x"3ed", x"3e3", x"3c8", x"39d", x"37f", x"368", x"365", x"373", x"38f", x"3af", x"3c9", x"3d3", 
			x"3cd", x"3c3", x"3ba", x"3b6", x"3b1", x"3b0", x"3aa", x"39c", x"38f", x"37d", x"37f", x"386", x"3a2", x"3c1", x"3d8", x"3dd", 
			x"3d1", x"3b3", x"399", x"381", x"37a", x"375", x"387", x"38b", x"38d", x"391", x"390", x"39f", x"3a7", x"3bf", x"3d1", x"3d5", 
			x"3ca", x"3b3", x"39d", x"38c", x"383", x"392", x"3a5", x"3bb", x"3e1", x"40b", x"418", x"432", x"416", x"3e9", x"3b3", x"379", 
			x"353", x"34b", x"34b", x"357", x"36d", x"384", x"390", x"3af", x"3b3", x"3b9", x"3b9", x"398", x"396", x"38c", x"39d", x"3a8", 
			x"3c7", x"3c0", x"3bc", x"3a7", x"397", x"393", x"3a7", x"3bc", x"3cf", x"3db", x"3c3", x"3a1", x"388", x"377", x"37e", x"393", 
			x"3b3", x"3c8", x"3db", x"3c2", x"3a8", x"392", x"37c", x"376", x"386", x"38e", x"3a8", x"3bd", x"3c1", x"3b3", x"3ab", x"3a8", 
			x"3ab", x"3b3", x"3b6", x"3c8", x"3be", x"3a7", x"391", x"381", x"37c", x"396", x"3b6", x"3d9", x"3ec", x"3df", x"3bf", x"398", 
			x"382", x"385", x"395", x"3ac", x"3c3", x"3be", x"3ad", x"395", x"385", x"389", x"392", x"3b4", x"3d8", x"3ef", x"3f6", x"3e9", 
			x"3df", x"3c6", x"3b6", x"39c", x"389", x"376", x"372", x"37a", x"396", x"3b4", x"3da", x"3ed", x"3f9", x"3e7", x"3d0", x"3b3", 
			x"39c", x"388", x"37b", x"374", x"374", x"37c", x"38b", x"3a2", x"3ab", x"3b4", x"3ab", x"3a5", x"3a5", x"3a6", x"39e", x"3a7", 
			x"39c", x"39c", x"399", x"397", x"3ab", x"3c3", x"3d3", x"3dd", x"3ce", x"3be", x"39e", x"393", x"390", x"39a", x"3aa", x"3b4", 
			x"3b7", x"3a4", x"395", x"387", x"387", x"391", x"3a6", x"3a7", x"3aa", x"3a6", x"3ab", x"3a8", x"3a9", x"3ad", x"3a5", x"397", 
			x"38f", x"38b", x"398", x"3b2", x"3e5", x"3f7", x"3fb", x"3de", x"3b0", x"380", x"364", x"35f", x"376", x"395", x"3ba", x"3d0", 
			x"3df", x"3d8", x"3c1", x"3b1", x"3a6", x"3a2", x"3a7", x"39d", x"39d", x"38b", x"383", x"37d", x"37c", x"38d", x"39c", x"3ae", 
			x"3bb", x"3b5", x"3b9", x"3ab", x"3b1", x"3ac", x"3b5", x"3ae", x"3a9", x"39f", x"399", x"3a0", x"3a0", x"3a8", x"3aa", x"3b2", 
			x"3be", x"3c9", x"3d4", x"3cf", x"3c1", x"3b1", x"3a2", x"39b", x"395", x"38b", x"38f", x"392", x"39d", x"3aa", x"3c1", x"3cb", 
			x"3ca", x"3b6", x"39f", x"389", x"38e", x"391", x"3a9", x"3d3", x"3f4", x"40a", x"406", x"3e3", x"3b4", x"393", x"383", x"380", 
			x"38d", x"39e", x"3b3", x"3bc", x"3c1", x"3cd", x"3cb", x"3d3", x"3cd", x"3c9", x"3b7", x"39b", x"387", x"379", x"371", x"372", 
			x"37d", x"38f", x"39f", x"3b1", x"3c8", x"3de", x"3e1", x"3d9", x"3c9", x"3aa", x"399", x"391", x"393", x"39f", x"3ab", x"3ab", 
			x"3b0", x"3af", x"3b9", x"3c7", x"3d2", x"3d4", x"3cb", x"3af", x"38b", x"375", x"36a", x"36f", x"37a", x"380", x"381", x"384", 
			x"37d", x"37b", x"384", x"38b", x"396", x"39d", x"3a3", x"39f", x"39c", x"38a", x"384", x"375", x"36e", x"372", x"388", x"39f", 
			x"3a1", x"3a4", x"399", x"392", x"387", x"378", x"383", x"38d", x"3a1", x"3ad", x"3a6", x"397", x"37f", x"37b", x"380", x"39f", 
			x"3b4", x"3ca", x"3b8", x"3b5", x"393", x"37e", x"384", x"390", x"39b", x"3b5", x"3d0", x"3ce", x"3c6", x"3b9", x"3b2", x"3b5", 
			x"3ae", x"3b0", x"3af", x"3a5", x"390", x"387", x"384", x"395", x"3aa", x"3b7", x"3ba", x"3a9", x"395", x"384", x"37f", x"379", 
			x"37f", x"389", x"397", x"3a5", x"39d", x"39a", x"38f", x"397", x"38a", x"389", x"39f", x"3a0", x"3ab", x"3ae", x"3a8", x"3af", 
			x"3bf", x"3bb", x"3b3", x"39f", x"38f", x"392", x"387", x"390", x"396", x"392", x"394", x"387", x"377", x"36d", x"377", x"38a", 
			x"3a9", x"3d7", x"3d9", x"3cc", x"3ab", x"388", x"373", x"36f", x"380", x"3a9", x"3c2", x"3e4", x"3e0", x"3c9", x"3b7", x"3ae", 
			x"3aa", x"3bb", x"3b8", x"3c7", x"3c3", x"3b2", x"3a2", x"394", x"38d", x"396", x"3b5", x"3c8", x"3d8", x"3cb", x"3ae", x"385", 
			x"36c", x"36b", x"36e", x"384", x"39f", x"3b6", x"3c4", x"3b8", x"3af", x"393", x"385", x"385", x"378", x"384", x"383", x"37d", 
			x"384", x"388", x"392", x"3aa", x"3c5", x"3e9", x"3e7", x"3cb", x"39d", x"37c", x"361", x"357", x"371", x"394", x"3b8", x"3c9", 
			x"3bf", x"3a6", x"38c", x"381", x"37b", x"389", x"392", x"394", x"38f", x"389", x"384", x"37f", x"38d", x"39e", x"3ac", x"3ba", 
			x"3c6", x"3cf", x"3d3", x"3df", x"3dc", x"3d1", x"3ca", x"3b5", x"3bd", x"3ad", x"3aa", x"3b8", x"3c2", x"3c7", x"3d1", x"3cc", 
			x"3d3", x"3cf", x"3d1", x"3c2", x"3bf", x"3ba", x"3b6", x"3ab", x"3af", x"3b8", x"3bf", x"3c7", x"3be", x"3b8", x"3ad", x"39d", 
			x"399", x"3b2", x"3be", x"3d3", x"3d0", x"3d3", x"3c1", x"3b3", x"3ab", x"3aa", x"3b8", x"3c3", x"3cd", x"3b0", x"3b3", x"38f", 
			x"391", x"3a2", x"3a1", x"3bf", x"3c8", x"3c9", x"3b5", x"3a3", x"3a6", x"39d", x"3ab", x"3a9", x"3c1", x"3b8", x"3cc", x"3b8", 
			x"3a2", x"3a0", x"398", x"3b7", x"3be", x"3e1", x"3f3", x"3f1", x"3f0", x"3f1", x"3e7", x"3d2", x"3d1", x"3ba", x"3b3", x"3ab", 
			x"3a6", x"3b8", x"3c3", x"3cf", x"3e0", x"3d2", x"3d8", x"3d7", x"3c4", x"3c7", x"3bc", x"3b5", x"3b7", x"3bd", x"3bf", x"3cf", 
			x"3c0", x"3c8", x"3bd", x"3b6", x"3b5", x"3c5", x"3db", x"3d8", x"3d7", x"3cf", x"3ba", x"3b0", x"3af", x"3b2", x"3c4", x"3cd", 
			x"3c0", x"3c5", x"3ad", x"3a5", x"39d", x"3a4", x"3b1", x"3ba", x"3c4", x"3c5", x"3c5", x"3b9", x"3ac", x"3aa", x"3af", x"3b8", 
			x"3c0", x"3b9", x"3bc", x"3c1", x"3af", x"3b0", x"3bb", x"3bd", x"3c5", x"3ba", x"3be", x"3ae", x"3ae", x"3a8", x"3b8", x"3c9", 
			x"3d9", x"3d5", x"3d8", x"3b3", x"3a3", x"39a", x"399", x"3a9", x"3b9", x"3cc", x"3cc", x"3b3", x"3a5", x"39a", x"3ad", x"3cf", 
			x"3e6", x"3ed", x"3da", x"3b1", x"399", x"38c", x"37e", x"39a", x"3ab", x"3c8", x"3d1", x"3d6", x"3dd", x"3de", x"3dd", x"3d0", 
			x"3c7", x"3ac", x"393", x"383", x"384", x"38a", x"3a0", x"3ca", x"3da", x"3dc", x"3ce", x"3b2", x"3a1", x"399", x"3a2", x"3b5", 
			x"3b6", x"3c7", x"3b8", x"3ac", x"398", x"39e", x"393", x"38f", x"3a0", x"3ad", x"3b7", x"3ce", x"3cd", x"3d4", x"3c0", x"3a6", 
			x"39a", x"398", x"39d", x"3ab", x"3bf", x"3be", x"3c2", x"3b1", x"3a1", x"39d", x"3a5", x"3a7", x"3b5", x"3a5", x"3a5", x"38e", 
			x"38d", x"391", x"39b", x"3c1", x"3d0", x"3d7", x"3c3", x"3ac", x"3a3", x"397", x"39a", x"3a1", x"39f", x"39b", x"398", x"3a5", 
			x"3aa", x"3bb", x"3cf", x"3dd", x"3d5", x"3b6", x"3a2", x"38b", x"383", x"383", x"38b", x"39b", x"3b0", x"3ad", x"3b6", x"3b9", 
			x"3a8", x"3af", x"39c", x"3a8", x"399", x"394", x"399", x"39a", x"3a9", x"3b2", x"3ad", x"3a0", x"397", x"38d", x"38d", x"39a", 
			x"3b6", x"3c3", x"3b8", x"3b9", x"3b2", x"397", x"38d", x"38c", x"38b", x"390", x"38b", x"391", x"3a4", x"3b1", x"3b9", x"3b8", 
			x"3b3", x"3a6", x"391", x"38f", x"380", x"38e", x"393", x"394", x"39a", x"3ac", x"3b4", x"3c3", x"3ba", x"3bf", x"3b3", x"3a0", 
			x"389", x"38e", x"392", x"39a", x"3ad", x"3b5", x"3b2", x"3b1", x"399", x"38e", x"390", x"39c", x"3a9", x"3a8", x"3a9", x"395", 
			x"387", x"378", x"38e", x"3a0", x"3bc", x"3d2", x"3d8", x"3c0", x"3a6", x"38f", x"38c", x"390", x"398", x"39f", x"3a4", x"3aa", 
			x"3b0", x"3b8", x"3b7", x"3bb", x"3ad", x"39f", x"39d", x"394", x"38c", x"397", x"395", x"395", x"395", x"390", x"390", x"397", 
			x"3ab", x"3bd", x"3cf", x"3c9", x"3b1", x"39a", x"389", x"383", x"380", x"388", x"397", x"39b", x"3a9", x"3b5", x"3bf", x"3cd", 
			x"3cc", x"3cc", x"3bb", x"39d", x"388", x"383", x"37c", x"38c", x"38f", x"3a9", x"3ac", x"3b3", x"3af", x"3a4", x"3a6", x"3a8", 
			x"39f", x"39a", x"394", x"38f", x"390", x"399", x"39f", x"3b3", x"3af", x"3a8", x"39f", x"393", x"39f", x"3ae", x"3b8", x"3b3", 
			x"3ab", x"3a5", x"3a1", x"3a4", x"3be", x"3ba", x"3be", x"3b0", x"397", x"386", x"383", x"393", x"3ab", x"3bb", x"3bf", x"3c4", 
			x"3ad", x"391", x"38e", x"38f", x"397", x"39f", x"3af", x"3b5", x"3af", x"3a0", x"391", x"38c", x"39e", x"398", x"3a7", x"3a3", 
			x"3a1", x"3ac", x"3a8", x"3b6", x"3b8", x"3bd", x"3b3", x"3a5", x"395", x"385", x"38f", x"391", x"39f", x"3ad", x"3b6", x"3b2", 
			x"3ab", x"3a2", x"3a7", x"3ac", x"3ac", x"3a7", x"391", x"381", x"37d", x"385", x"3a3", x"3b9", x"3c9", x"3c3", x"3bd", x"3af", 
			x"38c", x"385", x"37f", x"388", x"3a7", x"3b8", x"3c1", x"3c5", x"3c3", x"3af", x"3a7", x"3a0", x"3a4", x"3a8", x"3a4", x"3a2", 
			x"397", x"394", x"39c", x"399", x"3a8", x"3b5", x"3c3", x"3cd", x"3b9", x"3ab", x"396", x"37b", x"37b", x"381", x"396", x"3b9", 
			x"3d1", x"3e5", x"3d8", x"3c5", x"3a9", x"3eb", x"3bb", x"3bb", x"3d1", x"3f0", x"404", x"407", x"404", x"3f3", x"404", x"3fb", 
			x"3ef", x"3df", x"3f3", x"3f5", x"3e0", x"3cf", x"3ff", x"433", x"3e3", x"3a8", x"3a5", x"3ad", x"3c5", x"3cf", x"3d3", x"45a", 
			x"4cf", x"4cf", x"456", x"3ea", x"3cc", x"3cc", x"3da", x"42c", x"400", x"3f8", x"408", x"412", x"40e", x"3f0", x"3ee", x"409", 
			x"41c", x"40e", x"415", x"440", x"44a", x"43d", x"413", x"3f1", x"3e7", x"401", x"416", x"438", x"452", x"488", x"495", x"4e0", 
			x"4ad", x"463", x"435", x"42f", x"42f", x"43d", x"43c", x"431", x"41d", x"40d", x"40d", x"42b", x"44d", x"47d", x"471", x"475", 
			x"461", x"467", x"47b", x"497", x"4a5", x"495", x"480", x"457", x"44f", x"44a", x"465", x"47e", x"489", x"471", x"456", x"43e", 
			x"436", x"448", x"45c", x"46b", x"471", x"457", x"447", x"434", x"432", x"438", x"439", x"432", x"41a", x"406", x"3fb", x"3e5", 
			x"3d9", x"3d2", x"3c1", x"3a5", x"37d", x"35a", x"33b", x"324", x"316", x"300", x"2ea", x"2d6", x"2bd", x"2b9", x"2af", x"2ae", 
			x"2aa", x"2a7", x"29f", x"287", x"26b", x"255", x"244", x"23c", x"229", x"216", x"205", x"1f5", x"1d3", x"1b5", x"18f", x"16b", 
			x"143", x"129", x"120", x"124", x"133", x"15a", x"180", x"1b6", x"1de", x"1fa", x"208", x"235", x"260", x"290", x"2d2", x"32e", 
			x"364", x"390", x"3a6", x"3a1", x"3ca", x"3e3", x"3e7", x"3d9", x"3f4", x"429", x"434", x"40f", x"3fb", x"3d9", x"3f0", x"447", 
			x"497", x"4ca", x"4ee", x"4ee", x"4cb", x"486", x"469", x"458", x"419", x"37b", x"2fb", x"27b", x"211", x"1d6", x"1e4", x"1da", 
			x"1ce", x"1bc", x"1b5", x"1d6", x"1f1", x"249", x"2b0", x"2fa", x"351", x"44c", x"51c", x"5d2", x"5db", x"54a", x"4d7", x"3fc", 
			x"21c", x"0b7", x"015", x"11e", x"1e7", x"2a6", x"2ca", x"31f", x"3a8", x"407", x"481", x"4ca", x"430", x"2ef", x"29f", x"361", 
			x"38f", x"358", x"338", x"2bd", x"289", x"333", x"428", x"4e8", x"53d", x"580", x"5b0", x"5c1", x"5de", x"5ff", x"62f", x"64c", 
			x"65c", x"662", x"670", x"674", x"66e", x"667", x"658", x"621", x"5b9", x"57a", x"548", x"451", x"364", x"29a", x"2c5", x"35c", 
			x"2fa", x"267", x"22e", x"253", x"2af", x"31f", x"2aa", x"2d3", x"3df", x"581", x"5e8", x"574", x"4df", x"568", x"5ba", x"671", 
			x"6b1", x"6ca", x"69d", x"65f", x"61c", x"5ec", x"5c5", x"590", x"56f", x"5ae", x"67d", x"6e6", x"6c9", x"687", x"65b", x"663", 
			x"612", x"562", x"49b", x"439", x"440", x"3b2", x"2b9", x"2b8", x"2a5", x"2ac", x"236", x"233", x"297", x"343", x"449", x"517", 
			x"538", x"5aa", x"5b0", x"5e0", x"5e7", x"627", x"636", x"650", x"693", x"69f", x"668", x"68e", x"680", x"652", x"5e9", x"5ab", 
			x"587", x"578", x"549", x"51c", x"503", x"4ec", x"4ab", x"46d", x"458", x"460", x"464", x"459", x"478", x"501", x"599", x"5b5", 
			x"58e", x"532", x"4f8", x"4ee", x"50b", x"52a", x"564", x"589", x"5a8", x"56d", x"4b9", x"426", x"3bf", x"3c1", x"3f8", x"420", 
			x"46c", x"500", x"587", x"57b", x"56a", x"56d", x"5c2", x"5e6", x"593", x"544", x"52d", x"527", x"544", x"58f", x"5cc", x"66c", 
			x"70f", x"749", x"75b", x"757", x"730", x"6f8", x"6c4", x"6a4", x"696", x"67d", x"63f", x"5e8", x"599", x"556", x"52a", x"504", 
			x"4e4", x"4c5", x"49d", x"481", x"464", x"455", x"457", x"463", x"47f", x"49b", x"4c3", x"4e1", x"4c1", x"4a7", x"4b5", x"4ea", 
			x"53e", x"57c", x"5af", x"5d9", x"604", x"615", x"62c", x"64e", x"66e", x"683", x"68c", x"693", x"698", x"696", x"68b", x"674", 
			x"64e", x"645", x"638", x"633", x"625", x"5fc", x"5c9", x"598", x"56c", x"541", x"51c", x"4f9", x"4e5", x"4e3", x"4ea", x"502", 
			x"51a", x"517", x"4f0", x"4ca", x"4b0", x"4e5", x"55e", x"5ea", x"664", x"683", x"680", x"675", x"664", x"640", x"618", x"5e4", 
			x"5b1", x"583", x"57e", x"5c3", x"63d", x"6a9", x"6df", x"6f4", x"6f2", x"6cc", x"67d", x"627", x"5da", x"5a4", x"575", x"553", 
			x"53a", x"532", x"51f", x"502", x"4e5", x"4cf", x"4d6", x"4ee", x"511", x"559", x"5aa", x"5e5", x"610", x"624", x"618", x"5ee", 
			x"5b5", x"588", x"574", x"571", x"575", x"580", x"587", x"588", x"585", x"579", x"574", x"572", x"570", x"574", x"57a", x"584", 
			x"57f", x"573", x"563", x"558", x"546", x"53f", x"52f", x"528", x"520", x"519", x"50b", x"4fb", x"4f3", x"4ef", x"4f5", x"4f6", 
			x"4ef", x"4e6", x"4dd", x"4cf", x"4c6", x"4bf", x"4bf", x"4c6", x"4cb", x"4d8", x"4e3", x"4f1", x"4f9", x"4ff", x"512", x"51f", 
			x"538", x"54e", x"55b", x"56c", x"579", x"582", x"586", x"58f", x"593", x"590", x"588", x"575", x"554", x"52d", x"50b", x"4e3", 
			x"4ba", x"497", x"47a", x"464", x"451", x"449", x"43f", x"43f", x"43a", x"434", x"42a", x"41b", x"409", x"3f0", x"3de", x"3c9", 
			x"3c3", x"3bf", x"3c1", x"3c3", x"3cf", x"3d7", x"3e1", x"3e6", x"3ed", x"3ec", x"3e8", x"3e8", x"3df", x"3d7", x"3da", x"3e3", 
			x"3ec", x"3f8", x"406", x"410", x"41d", x"426", x"42f", x"438", x"43b", x"43d", x"43c", x"431", x"42f", x"42c", x"42c", x"431", 
			x"439", x"446", x"453", x"457", x"459", x"459", x"45c", x"463", x"469", x"473", x"47f", x"484", x"48d", x"48f", x"491", x"493", 
			x"49d", x"49d", x"49c", x"4a3", x"4a0", x"49e", x"49a", x"499", x"492", x"491", x"486", x"481", x"476", x"470", x"470", x"46e", 
			x"46c", x"467", x"464", x"464", x"460", x"45e", x"460", x"45e", x"461", x"468", x"467", x"46a", x"46a", x"46d", x"476", x"476", 
			x"474", x"475", x"471", x"46c", x"467", x"462", x"457", x"451", x"44b", x"445", x"43e", x"435", x"42a", x"428", x"423", x"41b", 
			x"416", x"413", x"40c", x"405", x"403", x"3fa", x"3f9", x"3f8", x"3ef", x"3ed", x"3e2", x"3e4", x"3db", x"3d3", x"3ce", x"3c9", 
			x"3c7", x"3c3", x"3c2", x"3c1", x"3c0", x"3c0", x"3c0", x"3c3", x"3c5", x"3c5", x"3c7", x"3c8", x"3c8", x"3c9", x"3c6", x"3ca", 
			x"3cb", x"3c9", x"3ca", x"3cf", x"3d0", x"3cb", x"3c5", x"3c7", x"3c4", x"3c7", x"3c6", x"3ca", x"3c5", x"3c2", x"3bd", x"3c3", 
			x"3c1", x"3be", x"3bd", x"3bf", x"3bd", x"3bf", x"3b7", x"3b8", x"3b3", x"3b2", x"3b1", x"3b1", x"3b4", x"3ae", x"3ab", x"3ac", 
			x"3aa", x"3a9", x"3ac", x"3af", x"3b0", x"3af", x"3b0", x"3b1", x"3ad", x"3ae", x"3aa", x"3aa", x"3a8", x"3a9", x"3a9", x"3a9", 
			x"3b0", x"3ad", x"3b3", x"3b0", x"3af", x"3b0", x"3af", x"3ae", x"3a9", x"3a9", x"3aa", x"3a9", x"3a7", x"3a4", x"39f", x"39a", 
			x"397", x"39a", x"394", x"38f", x"392", x"389", x"387", x"386", x"383", x"382", x"383", x"37d", x"378", x"376", x"372", x"376", 
			x"376", x"376", x"376", x"376", x"375", x"373", x"373", x"373", x"371", x"36d", x"373", x"36e", x"370", x"36e", x"373", x"36d", 
			x"370", x"36b", x"36d", x"36a", x"36e", x"370", x"369", x"369", x"365", x"363", x"35f", x"365", x"363", x"362", x"367", x"362", 
			x"360", x"35f", x"35e", x"35e", x"360", x"360", x"357", x"359", x"357", x"359", x"359", x"35a", x"35f", x"35e", x"35e", x"35d", 
			x"362", x"363", x"35d", x"35d", x"35d", x"35d", x"35c", x"35d", x"35e", x"360", x"35b", x"35d", x"35d", x"361", x"35b", x"35a", 
			x"35b", x"355", x"356", x"355", x"35b", x"35d", x"360", x"35f", x"35e", x"35e", x"35c", x"362", x"360", x"35e", x"363", x"361", 
			x"364", x"366", x"369", x"363", x"365", x"36d", x"36c", x"36d", x"36a", x"36e", x"36e", x"36d", x"367", x"36e", x"36e", x"36c", 
			x"36e", x"36c", x"372", x"373", x"372", x"372", x"36e", x"373", x"36d", x"36b", x"36b", x"36b", x"36a", x"36a", x"36c", x"36f", 
			x"374", x"374", x"373", x"372", x"36f", x"36f", x"36d", x"36b", x"36c", x"36e", x"368", x"36a", x"36b", x"366", x"364", x"36b", 
			x"366", x"367", x"369", x"369", x"366", x"367", x"368", x"36c", x"367", x"36d", x"36a", x"36a", x"36e", x"36b", x"36f", x"369", 
			x"36a", x"36b", x"36d", x"36c", x"36b", x"369", x"36c", x"369", x"36b", x"36b", x"366", x"364", x"369", x"367", x"369", x"36a", 
			x"36b", x"366", x"364", x"361", x"361", x"365", x"366", x"36a", x"36c", x"369", x"36c", x"36b", x"36b", x"366", x"366", x"363", 
			x"361", x"364", x"366", x"367", x"367", x"368", x"363", x"363", x"362", x"364", x"366", x"368", x"361", x"363", x"35f", x"364", 
			x"365", x"368", x"365", x"366", x"363", x"361", x"361", x"366", x"367", x"369", x"368", x"369", x"367", x"369", x"368", x"365", 
			x"368", x"368", x"369", x"36b", x"36a", x"36e", x"36c", x"369", x"368", x"36b", x"36b", x"36f", x"36d", x"36c", x"36e", x"36c", 
			x"36c", x"36d", x"36d", x"373", x"36f", x"36c", x"36c", x"36f", x"369", x"36f", x"36e", x"36d", x"370", x"371", x"371", x"373", 
			x"372", x"36f", x"375", x"372", x"370", x"374", x"372", x"372", x"372", x"36a", x"36e", x"375", x"378", x"37a", x"376", x"378", 
			x"374", x"372", x"374", x"372", x"374", x"374", x"376", x"371", x"371", x"36e", x"372", x"378", x"378", x"37c", x"37c", x"37e", 
			x"37c", x"37a", x"374", x"378", x"378", x"37b", x"37b", x"37d", x"37b", x"379", x"379", x"381", x"383", x"383", x"383", x"381", 
			x"382", x"380", x"37d", x"37d", x"380", x"388", x"388", x"38a", x"386", x"384", x"383", x"379", x"37b", x"383", x"382", x"37f", 
			x"386", x"37f", x"37f", x"382", x"380", x"37d", x"380", x"37e", x"37b", x"378", x"374", x"370", x"372", x"370", x"36f", x"377", 
			x"378", x"376", x"372", x"36f", x"36f", x"36b", x"36a", x"366", x"364", x"363", x"36b", x"367", x"362", x"362", x"361", x"35d", 
			x"361", x"365", x"365", x"35f", x"35b", x"35a", x"35c", x"360", x"35d", x"35d", x"363", x"35e", x"35e", x"35a", x"355", x"360", 
			x"35f", x"359", x"356", x"353", x"350", x"351", x"355", x"356", x"357", x"35e", x"35f", x"35e", x"35e", x"352", x"356", x"35e", 
			x"35a", x"35e", x"366", x"35e", x"362", x"35b", x"363", x"35c", x"363", x"360", x"368", x"36b", x"361", x"35f", x"35e", x"362", 
			x"35c", x"359", x"363", x"35c", x"367", x"35e", x"360", x"369", x"35e", x"368", x"363", x"367", x"363", x"365", x"35e", x"35b", 
			x"357", x"355", x"35f", x"35d", x"358", x"365", x"35b", x"356", x"354", x"354", x"35b", x"356", x"360", x"355", x"35b", x"360", 
			x"35b", x"35d", x"360", x"356", x"34e", x"35b", x"359", x"358", x"35b", x"359", x"358", x"357", x"359", x"355", x"358", x"357", 
			x"35b", x"35a", x"35d", x"34e", x"357", x"357", x"350", x"350", x"35b", x"34e", x"355", x"359", x"354", x"359", x"353", x"34d", 
			x"34e", x"350", x"34a", x"348", x"34a", x"34c", x"34c", x"34e", x"34c", x"348", x"345", x"346", x"344", x"345", x"341", x"33f", 
			x"33b", x"33b", x"33c", x"341", x"33e", x"342", x"341", x"341", x"341", x"33f", x"33e", x"33f", x"337", x"33b", x"341", x"33e", 
			x"345", x"346", x"34b", x"346", x"33f", x"33f", x"345", x"348", x"348", x"346", x"342", x"346", x"346", x"345", x"349", x"347", 
			x"34c", x"34b", x"349", x"344", x"345", x"347", x"348", x"348", x"34c", x"34c", x"354", x"353", x"354", x"359", x"351", x"34f", 
			x"352", x"351", x"34f", x"35c", x"359", x"359", x"35b", x"356", x"358", x"35b", x"359", x"35c", x"369", x"35f", x"356", x"356", 
			x"351", x"354", x"355", x"34e", x"34d", x"358", x"35a", x"35c", x"35f", x"35e", x"35f", x"352", x"354", x"355", x"34b", x"350", 
			x"355", x"361", x"361", x"35f", x"35b", x"365", x"35f", x"360", x"35f", x"35f", x"35b", x"359", x"357", x"357", x"364", x"36a", 
			x"36f", x"36f", x"376", x"36a", x"366", x"366", x"364", x"363", x"36d", x"36f", x"372", x"371", x"36b", x"368", x"36e", x"378", 
			x"371", x"372", x"36d", x"36f", x"371", x"366", x"365", x"36b", x"374", x"371", x"373", x"37b", x"37c", x"376", x"37b", x"371", 
			x"37a", x"36d", x"381", x"373", x"37e", x"375", x"375", x"373", x"376", x"375", x"374", x"37e", x"37e", x"37f", x"373", x"36f", 
			x"375", x"36f", x"36e", x"378", x"377", x"376", x"379", x"379", x"373", x"372", x"372", x"378", x"37c", x"376", x"378", x"376", 
			x"37a", x"378", x"37b", x"37a", x"383", x"38b", x"377", x"37b", x"37d", x"378", x"37f", x"375", x"379", x"380", x"380", x"38a", 
			x"383", x"382", x"384", x"37e", x"388", x"386", x"38e", x"38f", x"38a", x"392", x"38d", x"393", x"387", x"382", x"388", x"38d", 
			x"38e", x"38c", x"390", x"387", x"392", x"38c", x"38c", x"391", x"39d", x"39b", x"39e", x"39a", x"397", x"396", x"3a1", x"39c", 
			x"399", x"395", x"39b", x"396", x"396", x"398", x"399", x"39d", x"3a4", x"39c", x"398", x"397", x"394", x"394", x"398", x"39f", 
			x"395", x"399", x"393", x"395", x"395", x"39c", x"3a0", x"3a3", x"39b", x"398", x"394", x"396", x"38f", x"391", x"39a", x"39c", 
			x"398", x"395", x"395", x"392", x"393", x"38c", x"394", x"38f", x"38a", x"38a", x"383", x"387", x"380", x"388", x"388", x"38f", 
			x"388", x"397", x"38e", x"396", x"3a2", x"37f", x"386", x"38b", x"391", x"37d", x"383", x"382", x"393", x"382", x"381", x"388", 
			x"396", x"397", x"388", x"38a", x"389", x"387", x"37c", x"37a", x"387", x"385", x"38f", x"385", x"397", x"387", x"38b", x"38d", 
			x"384", x"383", x"383", x"37b", x"378", x"387", x"386", x"384", x"387", x"386", x"38b", x"38b", x"386", x"385", x"38d", x"389", 
			x"385", x"37f", x"389", x"388", x"384", x"38d", x"385", x"396", x"38a", x"38d", x"389", x"38c", x"386", x"38a", x"389", x"37e", 
			x"37e", x"37f", x"385", x"385", x"384", x"389", x"38b", x"38d", x"37f", x"381", x"384", x"37c", x"381", x"37a", x"380", x"377", 
			x"377", x"381", x"38a", x"38b", x"385", x"385", x"387", x"386", x"37c", x"37d", x"379", x"379", x"379", x"37f", x"386", x"38d", 
			x"389", x"386", x"38e", x"392", x"38c", x"386", x"389", x"38b", x"37e", x"37d", x"380", x"385", x"385", x"38f", x"389", x"383", 
			x"385", x"37a", x"384", x"37f", x"37f", x"381", x"385", x"382", x"382", x"37a", x"388", x"38a", x"392", x"38f", x"395", x"39a", 
			x"38f", x"390", x"381", x"388", x"37e", x"37e", x"382", x"38e", x"398", x"391", x"392", x"391", x"38e", x"38c", x"386", x"389", 
			x"390", x"38c", x"38b", x"382", x"380", x"38a", x"390", x"38e", x"398", x"392", x"390", x"383", x"384", x"37a", x"382", x"381", 
			x"38c", x"388", x"387", x"382", x"37e", x"37e", x"385", x"385", x"381", x"380", x"37b", x"37e", x"380", x"378", x"36e", x"376", 
			x"37c", x"37c", x"383", x"382", x"380", x"37a", x"37d", x"376", x"380", x"37c", x"375", x"374", x"379", x"370", x"379", x"380", 
			x"378", x"386", x"380", x"387", x"385", x"37f", x"383", x"37f", x"386", x"381", x"380", x"383", x"378", x"386", x"387", x"380", 
			x"38a", x"387", x"382", x"37f", x"380", x"37d", x"37c", x"381", x"383", x"37c", x"383", x"377", x"37c", x"381", x"38a", x"382", 
			x"384", x"382", x"37f", x"382", x"381", x"382", x"387", x"38d", x"38b", x"38b", x"38b", x"37f", x"38b", x"389", x"37e", x"383", 
			x"38b", x"382", x"380", x"37b", x"376", x"378", x"378", x"388", x"37e", x"384", x"393", x"38c", x"380", x"38c", x"378", x"37b", 
			x"37f", x"37e", x"37f", x"38c", x"38d", x"382", x"383", x"382", x"386", x"38d", x"392", x"389", x"38f", x"37d", x"384", x"384", 
			x"380", x"379", x"385", x"387", x"390", x"39d", x"395", x"399", x"38e", x"388", x"388", x"38a", x"38d", x"38c", x"38c", x"391", 
			x"391", x"399", x"393", x"38f", x"394", x"392", x"38b", x"396", x"38d", x"38e", x"382", x"391", x"388", x"393", x"399", x"39b", 
			x"397", x"396", x"398", x"39d", x"391", x"394", x"38d", x"38d", x"388", x"392", x"386", x"382", x"38f", x"388", x"384", x"388", 
			x"38b", x"381", x"38a", x"38b", x"388", x"391", x"391", x"38b", x"392", x"393", x"397", x"398", x"38f", x"399", x"38f", x"39b", 
			x"391", x"393", x"38e", x"38d", x"38e", x"38c", x"391", x"38f", x"396", x"384", x"38a", x"391", x"386", x"38d", x"387", x"37e", 
			x"38a", x"388", x"386", x"386", x"392", x"384", x"38c", x"38d", x"394", x"394", x"390", x"393", x"388", x"38a", x"384", x"391"
	);

	signal count : integer := 0;
	signal address : integer range 0 to ROM_LENGTH - 1 := 0;

begin

	dout <= DATA_ROM(address);

	process (clk, rst)
	begin
		if(rst = '1') then
			count <= 0;
			address <= 0;
		elsif(rising_edge(clk)) then
			count <= count + 1;
			
			if(count = 23) then
				if(address < ROM_LENGTH - 1) then
					address <= address + 1;
				else
					address <= 0;
				end if;
				
				count <= 0;
			end if;
		
		end if;
	end process;

end Behavioral;

